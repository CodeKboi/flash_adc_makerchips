* NGSPICE file created from priority_encoder.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

.subckt priority_encoder D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] O[0] O[1] O[2] O[3]
+ VGND VPWR clk
XTAP_TAPCELL_ROW_37_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput8 _18_/Q VGND VGND VPWR VPWR O[0] sky130_fd_sc_hd__buf_2
Xoutput10 _16_/Q VGND VGND VPWR VPWR O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 _17_/Q VGND VGND VPWR VPWR O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 _16_/CLK VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09_ _10_/C _10_/D VGND VGND VPWR VPWR _09_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08_ _11_/B VGND VGND VPWR VPWR _08_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_45_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpriority_encoder_11 VGND VGND VPWR VPWR priority_encoder_11/HI O[3] sky130_fd_sc_hd__conb_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 D[1] VGND VGND VPWR VPWR _13_/A2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 D[2] VGND VGND VPWR VPWR _11_/B sky130_fd_sc_hd__buf_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 D[3] VGND VGND VPWR VPWR _11_/A sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 D[4] VGND VGND VPWR VPWR _10_/D sky130_fd_sc_hd__buf_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 D[5] VGND VGND VPWR VPWR _10_/C sky130_fd_sc_hd__buf_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 D[6] VGND VGND VPWR VPWR _10_/B sky130_fd_sc_hd__buf_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 D[7] VGND VGND VPWR VPWR _10_/A sky130_fd_sc_hd__buf_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_62_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _18_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18_ _18_/CLK _18_/D VGND VGND VPWR VPWR _18_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17_ _18_/CLK _17_/D VGND VGND VPWR VPWR _17_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16_ _16_/CLK _16_/D VGND VGND VPWR VPWR _16_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _16_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15_ _10_/B _14_/X _10_/A VGND VGND VPWR VPWR _18_/D sky130_fd_sc_hd__o21bai_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14_ _10_/D _13_/Y _10_/C VGND VGND VPWR VPWR _14_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13_ _08_/Y _13_/A2 _11_/A VGND VGND VPWR VPWR _13_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12_ _09_/Y _11_/X _10_/A _10_/B VGND VGND VPWR VPWR _17_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11_ _11_/A _11_/B VGND VGND VPWR VPWR _11_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ _10_/A _10_/B _10_/C _10_/D VGND VGND VPWR VPWR _16_/D sky130_fd_sc_hd__or4_1
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends


magic
tech sky130A
magscale 1 2
timestamp 1730657462
<< nwell >>
rect 1066 2159 38862 37574
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< metal2 >>
rect 2594 39200 2650 40000
rect 7562 39200 7618 40000
rect 12530 39200 12586 40000
rect 17498 39200 17554 40000
rect 22466 39200 22522 40000
rect 27434 39200 27490 40000
rect 32402 39200 32458 40000
rect 37370 39200 37426 40000
rect 5078 0 5134 800
rect 15014 0 15070 800
rect 24950 0 25006 800
rect 34886 0 34942 800
<< obsm2 >>
rect 4214 39144 7506 39200
rect 7674 39144 12474 39200
rect 12642 39144 17442 39200
rect 17610 39144 22410 39200
rect 22578 39144 27378 39200
rect 27546 39144 32346 39200
rect 32514 39144 37314 39200
rect 37482 39144 37516 39200
rect 4214 856 37516 39144
rect 4214 800 5022 856
rect 5190 800 14958 856
rect 15126 800 24894 856
rect 25062 800 34830 856
rect 34998 800 37516 856
<< metal3 >>
rect 0 19864 800 19984
<< obsm3 >>
rect 800 20064 35246 37569
rect 880 19784 35246 20064
rect 800 2143 35246 19784
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 13675 19891 13741 27709
<< labels >>
rlabel metal2 s 2594 39200 2650 40000 6 D[0]
port 1 nsew signal input
rlabel metal2 s 7562 39200 7618 40000 6 D[1]
port 2 nsew signal input
rlabel metal2 s 12530 39200 12586 40000 6 D[2]
port 3 nsew signal input
rlabel metal2 s 17498 39200 17554 40000 6 D[3]
port 4 nsew signal input
rlabel metal2 s 22466 39200 22522 40000 6 D[4]
port 5 nsew signal input
rlabel metal2 s 27434 39200 27490 40000 6 D[5]
port 6 nsew signal input
rlabel metal2 s 32402 39200 32458 40000 6 D[6]
port 7 nsew signal input
rlabel metal2 s 37370 39200 37426 40000 6 D[7]
port 8 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 O[0]
port 9 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 O[1]
port 10 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 O[2]
port 11 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 O[3]
port 12 nsew signal output
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 13 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 14 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 14 nsew power bidirectional
rlabel metal3 s 0 19864 800 19984 6 clk
port 15 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 529970
string GDS_FILE /openlane/designs/encoder/runs/RUN_2024.11.03_18.10.17/results/signoff/priority_encoder.magic.gds
string GDS_START 106716
<< end >>


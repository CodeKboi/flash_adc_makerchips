magic
tech sky130A
magscale 1 2
timestamp 1730901471
<< checkpaint >>
rect -3932 -3932 13118 13932
<< viali >>
rect 5825 7497 5859 7531
rect 2053 7361 2087 7395
rect 3249 7361 3283 7395
rect 4629 7361 4663 7395
rect 5095 7361 5129 7395
rect 5273 7361 5307 7395
rect 5641 7361 5675 7395
rect 7021 7361 7055 7395
rect 8217 7361 8251 7395
rect 8493 7361 8527 7395
rect 2237 7157 2271 7191
rect 3433 7157 3467 7191
rect 4445 7157 4479 7191
rect 5273 7157 5307 7191
rect 6837 7157 6871 7191
rect 8033 7157 8067 7191
rect 8309 7157 8343 7191
rect 4445 6953 4479 6987
rect 6285 6953 6319 6987
rect 6193 6817 6227 6851
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 5927 6727 5961 6761
rect 6285 6749 6319 6783
rect 3893 6681 3927 6715
rect 6016 6681 6050 6715
rect 7113 6681 7147 6715
rect 3518 6613 3552 6647
rect 4261 6613 4295 6647
rect 5273 6613 5307 6647
rect 5365 6613 5399 6647
rect 6469 6613 6503 6647
rect 8033 6409 8067 6443
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 5457 6273 5491 6307
rect 6745 6273 6779 6307
rect 5181 6069 5215 6103
rect 6561 5661 6595 5695
rect 3617 5593 3651 5627
rect 4721 5593 4755 5627
rect 6806 5593 6840 5627
rect 2329 5525 2363 5559
rect 6009 5525 6043 5559
rect 7941 5525 7975 5559
rect 4068 5253 4102 5287
rect 3801 5117 3835 5151
rect 5181 4981 5215 5015
rect 5181 4573 5215 4607
rect 4936 4505 4970 4539
rect 3801 4437 3835 4471
rect 2053 2397 2087 2431
rect 5365 2397 5399 2431
rect 8217 2397 8251 2431
rect 1869 2261 1903 2295
rect 5181 2261 5215 2295
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 7642 8992 7664
rect 1104 7590 2882 7642
rect 2934 7590 2946 7642
rect 2998 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 4814 7642
rect 4866 7590 4878 7642
rect 4930 7590 4942 7642
rect 4994 7590 5006 7642
rect 5058 7590 5070 7642
rect 5122 7590 6746 7642
rect 6798 7590 6810 7642
rect 6862 7590 6874 7642
rect 6926 7590 6938 7642
rect 6990 7590 7002 7642
rect 7054 7590 8678 7642
rect 8730 7590 8742 7642
rect 8794 7590 8806 7642
rect 8858 7590 8870 7642
rect 8922 7590 8934 7642
rect 8986 7590 8992 7642
rect 1104 7568 8992 7590
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5276 7500 5825 7528
rect 5276 7404 5304 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 2038 7352 2044 7404
rect 2096 7352 2102 7404
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4396 7364 4629 7392
rect 4396 7352 4402 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 5074 7352 5080 7404
rect 5132 7401 5138 7404
rect 5132 7392 5141 7401
rect 5132 7364 5177 7392
rect 5132 7355 5141 7364
rect 5132 7352 5138 7355
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6696 7364 7021 7392
rect 6696 7352 6702 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7392 8539 7395
rect 9122 7392 9128 7404
rect 8527 7364 9128 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 3326 7188 3332 7200
rect 2271 7160 3332 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 3694 7188 3700 7200
rect 3467 7160 3700 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4304 7160 4445 7188
rect 4304 7148 4310 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4433 7151 4491 7157
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 5626 7188 5632 7200
rect 5307 7160 5632 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6236 7160 6837 7188
rect 6236 7148 6242 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 6972 7160 8033 7188
rect 6972 7148 6978 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8294 7148 8300 7200
rect 8352 7148 8358 7200
rect 1104 7098 8832 7120
rect 1104 7046 1916 7098
rect 1968 7046 1980 7098
rect 2032 7046 2044 7098
rect 2096 7046 2108 7098
rect 2160 7046 2172 7098
rect 2224 7046 3848 7098
rect 3900 7046 3912 7098
rect 3964 7046 3976 7098
rect 4028 7046 4040 7098
rect 4092 7046 4104 7098
rect 4156 7046 5780 7098
rect 5832 7046 5844 7098
rect 5896 7046 5908 7098
rect 5960 7046 5972 7098
rect 6024 7046 6036 7098
rect 6088 7046 7712 7098
rect 7764 7046 7776 7098
rect 7828 7046 7840 7098
rect 7892 7046 7904 7098
rect 7956 7046 7968 7098
rect 8020 7046 8832 7098
rect 1104 7024 8832 7046
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 3620 6956 4445 6984
rect 3620 6848 3648 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 4433 6947 4491 6953
rect 6273 6987 6331 6993
rect 6273 6953 6285 6987
rect 6319 6984 6331 6987
rect 6362 6984 6368 6996
rect 6319 6956 6368 6984
rect 6319 6953 6331 6956
rect 6273 6947 6331 6953
rect 6362 6944 6368 6956
rect 6420 6984 6426 6996
rect 6914 6984 6920 6996
rect 6420 6956 6920 6984
rect 6420 6944 6426 6956
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 5258 6916 5264 6928
rect 3752 6888 4384 6916
rect 3752 6876 3758 6888
rect 3436 6820 3648 6848
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 3436 6789 3464 6820
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3651 6752 4077 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 4065 6749 4077 6752
rect 4111 6780 4123 6783
rect 4246 6780 4252 6792
rect 4111 6752 4252 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4356 6789 4384 6888
rect 4632 6888 5264 6916
rect 4632 6789 4660 6888
rect 5258 6876 5264 6888
rect 5316 6876 5322 6928
rect 5368 6888 6224 6916
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3752 6684 3893 6712
rect 3752 6672 3758 6684
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 4816 6712 4844 6743
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5368 6780 5396 6888
rect 6196 6860 6224 6888
rect 5828 6820 6132 6848
rect 5828 6792 5856 6820
rect 5132 6752 5396 6780
rect 5537 6783 5595 6789
rect 5132 6740 5138 6752
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5552 6712 5580 6743
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 6104 6780 6132 6820
rect 6178 6808 6184 6860
rect 6236 6808 6242 6860
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5915 6761 5973 6767
rect 5915 6727 5927 6761
rect 5961 6727 5973 6761
rect 6104 6752 6285 6780
rect 6273 6749 6285 6752
rect 6319 6780 6331 6783
rect 8294 6780 8300 6792
rect 6319 6752 8300 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 5915 6724 5973 6727
rect 3881 6675 3939 6681
rect 4172 6684 4844 6712
rect 5092 6684 5580 6712
rect 3506 6647 3564 6653
rect 3506 6613 3518 6647
rect 3552 6644 3564 6647
rect 4172 6644 4200 6684
rect 3552 6616 4200 6644
rect 4249 6647 4307 6653
rect 3552 6613 3564 6616
rect 3506 6607 3564 6613
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 5092 6644 5120 6684
rect 5902 6672 5908 6724
rect 5960 6721 5973 6724
rect 5960 6672 5966 6721
rect 6004 6715 6062 6721
rect 6004 6681 6016 6715
rect 6050 6681 6062 6715
rect 6004 6675 6062 6681
rect 4295 6616 5120 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 5224 6616 5273 6644
rect 5224 6604 5230 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6012 6644 6040 6675
rect 7098 6672 7104 6724
rect 7156 6672 7162 6724
rect 5500 6616 6040 6644
rect 5500 6604 5506 6616
rect 6454 6604 6460 6656
rect 6512 6604 6518 6656
rect 1104 6554 8992 6576
rect 1104 6502 2882 6554
rect 2934 6502 2946 6554
rect 2998 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 4814 6554
rect 4866 6502 4878 6554
rect 4930 6502 4942 6554
rect 4994 6502 5006 6554
rect 5058 6502 5070 6554
rect 5122 6502 6746 6554
rect 6798 6502 6810 6554
rect 6862 6502 6874 6554
rect 6926 6502 6938 6554
rect 6990 6502 7002 6554
rect 7054 6502 8678 6554
rect 8730 6502 8742 6554
rect 8794 6502 8806 6554
rect 8858 6502 8870 6554
rect 8922 6502 8934 6554
rect 8986 6502 8992 6554
rect 1104 6480 8992 6502
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7156 6412 8033 6440
rect 7156 6400 7162 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 5902 6372 5908 6384
rect 5000 6344 5908 6372
rect 5000 6313 5028 6344
rect 5902 6332 5908 6344
rect 5960 6372 5966 6384
rect 6362 6372 6368 6384
rect 5960 6344 6368 6372
rect 5960 6332 5966 6344
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5810 6304 5816 6316
rect 5491 6276 5816 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6696 6276 6745 6304
rect 6696 6264 6702 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 1104 6010 8832 6032
rect 1104 5958 1916 6010
rect 1968 5958 1980 6010
rect 2032 5958 2044 6010
rect 2096 5958 2108 6010
rect 2160 5958 2172 6010
rect 2224 5958 3848 6010
rect 3900 5958 3912 6010
rect 3964 5958 3976 6010
rect 4028 5958 4040 6010
rect 4092 5958 4104 6010
rect 4156 5958 5780 6010
rect 5832 5958 5844 6010
rect 5896 5958 5908 6010
rect 5960 5958 5972 6010
rect 6024 5958 6036 6010
rect 6088 5958 7712 6010
rect 7764 5958 7776 6010
rect 7828 5958 7840 6010
rect 7892 5958 7904 6010
rect 7956 5958 7968 6010
rect 8020 5958 8832 6010
rect 1104 5936 8832 5958
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 7098 5692 7104 5704
rect 6595 5664 7104 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 3605 5627 3663 5633
rect 3605 5593 3617 5627
rect 3651 5624 3663 5627
rect 3651 5596 4108 5624
rect 3651 5593 3663 5596
rect 3605 5587 3663 5593
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 3694 5556 3700 5568
rect 2363 5528 3700 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 4080 5556 4108 5596
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4709 5627 4767 5633
rect 4709 5624 4721 5627
rect 4212 5596 4721 5624
rect 4212 5584 4218 5596
rect 4709 5593 4721 5596
rect 4755 5593 4767 5627
rect 4709 5587 4767 5593
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 6794 5627 6852 5633
rect 6794 5624 6806 5627
rect 6512 5596 6806 5624
rect 6512 5584 6518 5596
rect 6794 5593 6806 5596
rect 6840 5593 6852 5627
rect 6794 5587 6852 5593
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 4080 5528 6009 5556
rect 5997 5525 6009 5528
rect 6043 5556 6055 5559
rect 6638 5556 6644 5568
rect 6043 5528 6644 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 8202 5556 8208 5568
rect 7975 5528 8208 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 1104 5466 8992 5488
rect 1104 5414 2882 5466
rect 2934 5414 2946 5466
rect 2998 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 4814 5466
rect 4866 5414 4878 5466
rect 4930 5414 4942 5466
rect 4994 5414 5006 5466
rect 5058 5414 5070 5466
rect 5122 5414 6746 5466
rect 6798 5414 6810 5466
rect 6862 5414 6874 5466
rect 6926 5414 6938 5466
rect 6990 5414 7002 5466
rect 7054 5414 8678 5466
rect 8730 5414 8742 5466
rect 8794 5414 8806 5466
rect 8858 5414 8870 5466
rect 8922 5414 8934 5466
rect 8986 5414 8992 5466
rect 1104 5392 8992 5414
rect 4056 5287 4114 5293
rect 4056 5253 4068 5287
rect 4102 5284 4114 5287
rect 5350 5284 5356 5296
rect 4102 5256 5356 5284
rect 4102 5253 4114 5256
rect 4056 5247 4114 5253
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3752 5120 3801 5148
rect 3752 5108 3758 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 5012 5227 5015
rect 5350 5012 5356 5024
rect 5215 4984 5356 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 1104 4922 8832 4944
rect 1104 4870 1916 4922
rect 1968 4870 1980 4922
rect 2032 4870 2044 4922
rect 2096 4870 2108 4922
rect 2160 4870 2172 4922
rect 2224 4870 3848 4922
rect 3900 4870 3912 4922
rect 3964 4870 3976 4922
rect 4028 4870 4040 4922
rect 4092 4870 4104 4922
rect 4156 4870 5780 4922
rect 5832 4870 5844 4922
rect 5896 4870 5908 4922
rect 5960 4870 5972 4922
rect 6024 4870 6036 4922
rect 6088 4870 7712 4922
rect 7764 4870 7776 4922
rect 7828 4870 7840 4922
rect 7892 4870 7904 4922
rect 7956 4870 7968 4922
rect 8020 4870 8832 4922
rect 1104 4848 8832 4870
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 3752 4576 5181 4604
rect 3752 4564 3758 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 4924 4539 4982 4545
rect 4924 4505 4936 4539
rect 4970 4536 4982 4539
rect 5074 4536 5080 4548
rect 4970 4508 5080 4536
rect 4970 4505 4982 4508
rect 4924 4499 4982 4505
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 2832 4440 3801 4468
rect 2832 4428 2838 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 1104 4378 8992 4400
rect 1104 4326 2882 4378
rect 2934 4326 2946 4378
rect 2998 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 4814 4378
rect 4866 4326 4878 4378
rect 4930 4326 4942 4378
rect 4994 4326 5006 4378
rect 5058 4326 5070 4378
rect 5122 4326 6746 4378
rect 6798 4326 6810 4378
rect 6862 4326 6874 4378
rect 6926 4326 6938 4378
rect 6990 4326 7002 4378
rect 7054 4326 8678 4378
rect 8730 4326 8742 4378
rect 8794 4326 8806 4378
rect 8858 4326 8870 4378
rect 8922 4326 8934 4378
rect 8986 4326 8992 4378
rect 1104 4304 8992 4326
rect 1104 3834 8832 3856
rect 1104 3782 1916 3834
rect 1968 3782 1980 3834
rect 2032 3782 2044 3834
rect 2096 3782 2108 3834
rect 2160 3782 2172 3834
rect 2224 3782 3848 3834
rect 3900 3782 3912 3834
rect 3964 3782 3976 3834
rect 4028 3782 4040 3834
rect 4092 3782 4104 3834
rect 4156 3782 5780 3834
rect 5832 3782 5844 3834
rect 5896 3782 5908 3834
rect 5960 3782 5972 3834
rect 6024 3782 6036 3834
rect 6088 3782 7712 3834
rect 7764 3782 7776 3834
rect 7828 3782 7840 3834
rect 7892 3782 7904 3834
rect 7956 3782 7968 3834
rect 8020 3782 8832 3834
rect 1104 3760 8832 3782
rect 1104 3290 8992 3312
rect 1104 3238 2882 3290
rect 2934 3238 2946 3290
rect 2998 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 4814 3290
rect 4866 3238 4878 3290
rect 4930 3238 4942 3290
rect 4994 3238 5006 3290
rect 5058 3238 5070 3290
rect 5122 3238 6746 3290
rect 6798 3238 6810 3290
rect 6862 3238 6874 3290
rect 6926 3238 6938 3290
rect 6990 3238 7002 3290
rect 7054 3238 8678 3290
rect 8730 3238 8742 3290
rect 8794 3238 8806 3290
rect 8858 3238 8870 3290
rect 8922 3238 8934 3290
rect 8986 3238 8992 3290
rect 1104 3216 8992 3238
rect 1104 2746 8832 2768
rect 1104 2694 1916 2746
rect 1968 2694 1980 2746
rect 2032 2694 2044 2746
rect 2096 2694 2108 2746
rect 2160 2694 2172 2746
rect 2224 2694 3848 2746
rect 3900 2694 3912 2746
rect 3964 2694 3976 2746
rect 4028 2694 4040 2746
rect 4092 2694 4104 2746
rect 4156 2694 5780 2746
rect 5832 2694 5844 2746
rect 5896 2694 5908 2746
rect 5960 2694 5972 2746
rect 6024 2694 6036 2746
rect 6088 2694 7712 2746
rect 7764 2694 7776 2746
rect 7828 2694 7840 2746
rect 7892 2694 7904 2746
rect 7956 2694 7968 2746
rect 8020 2694 8832 2746
rect 1104 2672 8832 2694
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2774 2428 2780 2440
rect 2087 2400 2780 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 1728 2264 1869 2292
rect 1728 2252 1734 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 5166 2252 5172 2304
rect 5224 2252 5230 2304
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8389 2295 8447 2301
rect 8389 2292 8401 2295
rect 8352 2264 8401 2292
rect 8352 2252 8358 2264
rect 8389 2261 8401 2264
rect 8435 2261 8447 2295
rect 8389 2255 8447 2261
rect 1104 2202 8992 2224
rect 1104 2150 2882 2202
rect 2934 2150 2946 2202
rect 2998 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 4814 2202
rect 4866 2150 4878 2202
rect 4930 2150 4942 2202
rect 4994 2150 5006 2202
rect 5058 2150 5070 2202
rect 5122 2150 6746 2202
rect 6798 2150 6810 2202
rect 6862 2150 6874 2202
rect 6926 2150 6938 2202
rect 6990 2150 7002 2202
rect 7054 2150 8678 2202
rect 8730 2150 8742 2202
rect 8794 2150 8806 2202
rect 8858 2150 8870 2202
rect 8922 2150 8934 2202
rect 8986 2150 8992 2202
rect 1104 2128 8992 2150
<< via1 >>
rect 2882 7590 2934 7642
rect 2946 7590 2998 7642
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 4814 7590 4866 7642
rect 4878 7590 4930 7642
rect 4942 7590 4994 7642
rect 5006 7590 5058 7642
rect 5070 7590 5122 7642
rect 6746 7590 6798 7642
rect 6810 7590 6862 7642
rect 6874 7590 6926 7642
rect 6938 7590 6990 7642
rect 7002 7590 7054 7642
rect 8678 7590 8730 7642
rect 8742 7590 8794 7642
rect 8806 7590 8858 7642
rect 8870 7590 8922 7642
rect 8934 7590 8986 7642
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 4344 7352 4396 7404
rect 5080 7395 5132 7404
rect 5080 7361 5095 7395
rect 5095 7361 5129 7395
rect 5129 7361 5132 7395
rect 5080 7352 5132 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5540 7352 5592 7404
rect 6644 7352 6696 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 9128 7352 9180 7404
rect 3332 7148 3384 7200
rect 3700 7148 3752 7200
rect 4252 7148 4304 7200
rect 5632 7148 5684 7200
rect 6184 7148 6236 7200
rect 6920 7148 6972 7200
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 1916 7046 1968 7098
rect 1980 7046 2032 7098
rect 2044 7046 2096 7098
rect 2108 7046 2160 7098
rect 2172 7046 2224 7098
rect 3848 7046 3900 7098
rect 3912 7046 3964 7098
rect 3976 7046 4028 7098
rect 4040 7046 4092 7098
rect 4104 7046 4156 7098
rect 5780 7046 5832 7098
rect 5844 7046 5896 7098
rect 5908 7046 5960 7098
rect 5972 7046 6024 7098
rect 6036 7046 6088 7098
rect 7712 7046 7764 7098
rect 7776 7046 7828 7098
rect 7840 7046 7892 7098
rect 7904 7046 7956 7098
rect 7968 7046 8020 7098
rect 6368 6944 6420 6996
rect 6920 6944 6972 6996
rect 3700 6876 3752 6928
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4252 6740 4304 6792
rect 5264 6876 5316 6928
rect 3700 6672 3752 6724
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 8300 6740 8352 6792
rect 5908 6672 5960 6724
rect 5172 6604 5224 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 5448 6604 5500 6656
rect 7104 6715 7156 6724
rect 7104 6681 7113 6715
rect 7113 6681 7147 6715
rect 7147 6681 7156 6715
rect 7104 6672 7156 6681
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 2882 6502 2934 6554
rect 2946 6502 2998 6554
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 4814 6502 4866 6554
rect 4878 6502 4930 6554
rect 4942 6502 4994 6554
rect 5006 6502 5058 6554
rect 5070 6502 5122 6554
rect 6746 6502 6798 6554
rect 6810 6502 6862 6554
rect 6874 6502 6926 6554
rect 6938 6502 6990 6554
rect 7002 6502 7054 6554
rect 8678 6502 8730 6554
rect 8742 6502 8794 6554
rect 8806 6502 8858 6554
rect 8870 6502 8922 6554
rect 8934 6502 8986 6554
rect 7104 6400 7156 6452
rect 5908 6332 5960 6384
rect 6368 6332 6420 6384
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5816 6264 5868 6316
rect 6644 6264 6696 6316
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 1916 5958 1968 6010
rect 1980 5958 2032 6010
rect 2044 5958 2096 6010
rect 2108 5958 2160 6010
rect 2172 5958 2224 6010
rect 3848 5958 3900 6010
rect 3912 5958 3964 6010
rect 3976 5958 4028 6010
rect 4040 5958 4092 6010
rect 4104 5958 4156 6010
rect 5780 5958 5832 6010
rect 5844 5958 5896 6010
rect 5908 5958 5960 6010
rect 5972 5958 6024 6010
rect 6036 5958 6088 6010
rect 7712 5958 7764 6010
rect 7776 5958 7828 6010
rect 7840 5958 7892 6010
rect 7904 5958 7956 6010
rect 7968 5958 8020 6010
rect 7104 5652 7156 5704
rect 3700 5516 3752 5568
rect 4160 5584 4212 5636
rect 6460 5584 6512 5636
rect 6644 5516 6696 5568
rect 8208 5516 8260 5568
rect 2882 5414 2934 5466
rect 2946 5414 2998 5466
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 4814 5414 4866 5466
rect 4878 5414 4930 5466
rect 4942 5414 4994 5466
rect 5006 5414 5058 5466
rect 5070 5414 5122 5466
rect 6746 5414 6798 5466
rect 6810 5414 6862 5466
rect 6874 5414 6926 5466
rect 6938 5414 6990 5466
rect 7002 5414 7054 5466
rect 8678 5414 8730 5466
rect 8742 5414 8794 5466
rect 8806 5414 8858 5466
rect 8870 5414 8922 5466
rect 8934 5414 8986 5466
rect 5356 5244 5408 5296
rect 3700 5108 3752 5160
rect 5356 4972 5408 5024
rect 1916 4870 1968 4922
rect 1980 4870 2032 4922
rect 2044 4870 2096 4922
rect 2108 4870 2160 4922
rect 2172 4870 2224 4922
rect 3848 4870 3900 4922
rect 3912 4870 3964 4922
rect 3976 4870 4028 4922
rect 4040 4870 4092 4922
rect 4104 4870 4156 4922
rect 5780 4870 5832 4922
rect 5844 4870 5896 4922
rect 5908 4870 5960 4922
rect 5972 4870 6024 4922
rect 6036 4870 6088 4922
rect 7712 4870 7764 4922
rect 7776 4870 7828 4922
rect 7840 4870 7892 4922
rect 7904 4870 7956 4922
rect 7968 4870 8020 4922
rect 3700 4564 3752 4616
rect 5080 4496 5132 4548
rect 2780 4428 2832 4480
rect 2882 4326 2934 4378
rect 2946 4326 2998 4378
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 4814 4326 4866 4378
rect 4878 4326 4930 4378
rect 4942 4326 4994 4378
rect 5006 4326 5058 4378
rect 5070 4326 5122 4378
rect 6746 4326 6798 4378
rect 6810 4326 6862 4378
rect 6874 4326 6926 4378
rect 6938 4326 6990 4378
rect 7002 4326 7054 4378
rect 8678 4326 8730 4378
rect 8742 4326 8794 4378
rect 8806 4326 8858 4378
rect 8870 4326 8922 4378
rect 8934 4326 8986 4378
rect 1916 3782 1968 3834
rect 1980 3782 2032 3834
rect 2044 3782 2096 3834
rect 2108 3782 2160 3834
rect 2172 3782 2224 3834
rect 3848 3782 3900 3834
rect 3912 3782 3964 3834
rect 3976 3782 4028 3834
rect 4040 3782 4092 3834
rect 4104 3782 4156 3834
rect 5780 3782 5832 3834
rect 5844 3782 5896 3834
rect 5908 3782 5960 3834
rect 5972 3782 6024 3834
rect 6036 3782 6088 3834
rect 7712 3782 7764 3834
rect 7776 3782 7828 3834
rect 7840 3782 7892 3834
rect 7904 3782 7956 3834
rect 7968 3782 8020 3834
rect 2882 3238 2934 3290
rect 2946 3238 2998 3290
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 4814 3238 4866 3290
rect 4878 3238 4930 3290
rect 4942 3238 4994 3290
rect 5006 3238 5058 3290
rect 5070 3238 5122 3290
rect 6746 3238 6798 3290
rect 6810 3238 6862 3290
rect 6874 3238 6926 3290
rect 6938 3238 6990 3290
rect 7002 3238 7054 3290
rect 8678 3238 8730 3290
rect 8742 3238 8794 3290
rect 8806 3238 8858 3290
rect 8870 3238 8922 3290
rect 8934 3238 8986 3290
rect 1916 2694 1968 2746
rect 1980 2694 2032 2746
rect 2044 2694 2096 2746
rect 2108 2694 2160 2746
rect 2172 2694 2224 2746
rect 3848 2694 3900 2746
rect 3912 2694 3964 2746
rect 3976 2694 4028 2746
rect 4040 2694 4092 2746
rect 4104 2694 4156 2746
rect 5780 2694 5832 2746
rect 5844 2694 5896 2746
rect 5908 2694 5960 2746
rect 5972 2694 6024 2746
rect 6036 2694 6088 2746
rect 7712 2694 7764 2746
rect 7776 2694 7828 2746
rect 7840 2694 7892 2746
rect 7904 2694 7956 2746
rect 7968 2694 8020 2746
rect 2780 2388 2832 2440
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 1676 2252 1728 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 8300 2252 8352 2304
rect 2882 2150 2934 2202
rect 2946 2150 2998 2202
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 4814 2150 4866 2202
rect 4878 2150 4930 2202
rect 4942 2150 4994 2202
rect 5006 2150 5058 2202
rect 5070 2150 5122 2202
rect 6746 2150 6798 2202
rect 6810 2150 6862 2202
rect 6874 2150 6926 2202
rect 6938 2150 6990 2202
rect 7002 2150 7054 2202
rect 8678 2150 8730 2202
rect 8742 2150 8794 2202
rect 8806 2150 8858 2202
rect 8870 2150 8922 2202
rect 8934 2150 8986 2202
<< metal2 >>
rect 754 9200 810 10000
rect 1950 9330 2006 10000
rect 3146 9330 3202 10000
rect 1950 9302 2084 9330
rect 1950 9200 2006 9302
rect 2056 7410 2084 9302
rect 3146 9302 3280 9330
rect 3146 9200 3202 9302
rect 2882 7644 3190 7653
rect 2882 7642 2888 7644
rect 2944 7642 2968 7644
rect 3024 7642 3048 7644
rect 3104 7642 3128 7644
rect 3184 7642 3190 7644
rect 2944 7590 2946 7642
rect 3126 7590 3128 7642
rect 2882 7588 2888 7590
rect 2944 7588 2968 7590
rect 3024 7588 3048 7590
rect 3104 7588 3128 7590
rect 3184 7588 3190 7590
rect 2882 7579 3190 7588
rect 3252 7410 3280 9302
rect 4342 9200 4398 10000
rect 5538 9200 5594 10000
rect 6734 9200 6790 10000
rect 7930 9330 7986 10000
rect 7930 9302 8248 9330
rect 7930 9200 7986 9302
rect 4356 7410 4384 9200
rect 4814 7644 5122 7653
rect 4814 7642 4820 7644
rect 4876 7642 4900 7644
rect 4956 7642 4980 7644
rect 5036 7642 5060 7644
rect 5116 7642 5122 7644
rect 4876 7590 4878 7642
rect 5058 7590 5060 7642
rect 4814 7588 4820 7590
rect 4876 7588 4900 7590
rect 4956 7588 4980 7590
rect 5036 7588 5060 7590
rect 5116 7588 5122 7590
rect 4814 7579 5122 7588
rect 5552 7410 5580 9200
rect 6748 7834 6776 9200
rect 6656 7806 6776 7834
rect 6656 7410 6684 7806
rect 6746 7644 7054 7653
rect 6746 7642 6752 7644
rect 6808 7642 6832 7644
rect 6888 7642 6912 7644
rect 6968 7642 6992 7644
rect 7048 7642 7054 7644
rect 6808 7590 6810 7642
rect 6990 7590 6992 7642
rect 6746 7588 6752 7590
rect 6808 7588 6832 7590
rect 6888 7588 6912 7590
rect 6968 7588 6992 7590
rect 7048 7588 7054 7590
rect 6746 7579 7054 7588
rect 8220 7410 8248 9302
rect 9126 9200 9182 10000
rect 8678 7644 8986 7653
rect 8678 7642 8684 7644
rect 8740 7642 8764 7644
rect 8820 7642 8844 7644
rect 8900 7642 8924 7644
rect 8980 7642 8986 7644
rect 8740 7590 8742 7642
rect 8922 7590 8924 7642
rect 8678 7588 8684 7590
rect 8740 7588 8764 7590
rect 8820 7588 8844 7590
rect 8900 7588 8924 7590
rect 8980 7588 8986 7590
rect 8678 7579 8986 7588
rect 9140 7410 9168 9200
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 1916 7100 2224 7109
rect 1916 7098 1922 7100
rect 1978 7098 2002 7100
rect 2058 7098 2082 7100
rect 2138 7098 2162 7100
rect 2218 7098 2224 7100
rect 1978 7046 1980 7098
rect 2160 7046 2162 7098
rect 1916 7044 1922 7046
rect 1978 7044 2002 7046
rect 2058 7044 2082 7046
rect 2138 7044 2162 7046
rect 2218 7044 2224 7046
rect 1916 7035 2224 7044
rect 3344 6798 3372 7142
rect 3712 6934 3740 7142
rect 3848 7100 4156 7109
rect 3848 7098 3854 7100
rect 3910 7098 3934 7100
rect 3990 7098 4014 7100
rect 4070 7098 4094 7100
rect 4150 7098 4156 7100
rect 3910 7046 3912 7098
rect 4092 7046 4094 7098
rect 3848 7044 3854 7046
rect 3910 7044 3934 7046
rect 3990 7044 4014 7046
rect 4070 7044 4094 7046
rect 4150 7044 4156 7046
rect 3848 7035 4156 7044
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3712 6730 3740 6870
rect 4264 6798 4292 7142
rect 5092 6798 5120 7346
rect 5276 6934 5304 7346
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 5264 6928 5316 6934
rect 5316 6888 5488 6916
rect 5264 6870 5316 6876
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 5460 6662 5488 6888
rect 5644 6798 5672 7142
rect 5780 7100 6088 7109
rect 5780 7098 5786 7100
rect 5842 7098 5866 7100
rect 5922 7098 5946 7100
rect 6002 7098 6026 7100
rect 6082 7098 6088 7100
rect 5842 7046 5844 7098
rect 6024 7046 6026 7098
rect 5780 7044 5786 7046
rect 5842 7044 5866 7046
rect 5922 7044 5946 7046
rect 6002 7044 6026 7046
rect 6082 7044 6088 7046
rect 5780 7035 6088 7044
rect 6196 6866 6224 7142
rect 6932 7002 6960 7142
rect 7712 7100 8020 7109
rect 7712 7098 7718 7100
rect 7774 7098 7798 7100
rect 7854 7098 7878 7100
rect 7934 7098 7958 7100
rect 8014 7098 8020 7100
rect 7774 7046 7776 7098
rect 7956 7046 7958 7098
rect 7712 7044 7718 7046
rect 7774 7044 7798 7046
rect 7854 7044 7878 7046
rect 7934 7044 7958 7046
rect 8014 7044 8020 7046
rect 7712 7035 8020 7044
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 2882 6556 3190 6565
rect 2882 6554 2888 6556
rect 2944 6554 2968 6556
rect 3024 6554 3048 6556
rect 3104 6554 3128 6556
rect 3184 6554 3190 6556
rect 2944 6502 2946 6554
rect 3126 6502 3128 6554
rect 2882 6500 2888 6502
rect 2944 6500 2968 6502
rect 3024 6500 3048 6502
rect 3104 6500 3128 6502
rect 3184 6500 3190 6502
rect 2882 6491 3190 6500
rect 4814 6556 5122 6565
rect 4814 6554 4820 6556
rect 4876 6554 4900 6556
rect 4956 6554 4980 6556
rect 5036 6554 5060 6556
rect 5116 6554 5122 6556
rect 4876 6502 4878 6554
rect 5058 6502 5060 6554
rect 4814 6500 4820 6502
rect 4876 6500 4900 6502
rect 4956 6500 4980 6502
rect 5036 6500 5060 6502
rect 5116 6500 5122 6502
rect 4814 6491 5122 6500
rect 5184 6322 5212 6598
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 1916 6012 2224 6021
rect 1916 6010 1922 6012
rect 1978 6010 2002 6012
rect 2058 6010 2082 6012
rect 2138 6010 2162 6012
rect 2218 6010 2224 6012
rect 1978 5958 1980 6010
rect 2160 5958 2162 6010
rect 1916 5956 1922 5958
rect 1978 5956 2002 5958
rect 2058 5956 2082 5958
rect 2138 5956 2162 5958
rect 2218 5956 2224 5958
rect 1916 5947 2224 5956
rect 3848 6012 4156 6021
rect 3848 6010 3854 6012
rect 3910 6010 3934 6012
rect 3990 6010 4014 6012
rect 4070 6010 4094 6012
rect 4150 6010 4156 6012
rect 3910 5958 3912 6010
rect 4092 5958 4094 6010
rect 3848 5956 3854 5958
rect 3910 5956 3934 5958
rect 3990 5956 4014 5958
rect 4070 5956 4094 5958
rect 4150 5956 4156 5958
rect 3848 5947 4156 5956
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 2882 5468 3190 5477
rect 2882 5466 2888 5468
rect 2944 5466 2968 5468
rect 3024 5466 3048 5468
rect 3104 5466 3128 5468
rect 3184 5466 3190 5468
rect 2944 5414 2946 5466
rect 3126 5414 3128 5466
rect 2882 5412 2888 5414
rect 2944 5412 2968 5414
rect 3024 5412 3048 5414
rect 3104 5412 3128 5414
rect 3184 5412 3190 5414
rect 2882 5403 3190 5412
rect 3712 5166 3740 5510
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 4066 5128 4122 5137
rect 1916 4924 2224 4933
rect 1916 4922 1922 4924
rect 1978 4922 2002 4924
rect 2058 4922 2082 4924
rect 2138 4922 2162 4924
rect 2218 4922 2224 4924
rect 1978 4870 1980 4922
rect 2160 4870 2162 4922
rect 1916 4868 1922 4870
rect 1978 4868 2002 4870
rect 2058 4868 2082 4870
rect 2138 4868 2162 4870
rect 2218 4868 2224 4870
rect 1916 4859 2224 4868
rect 3712 4622 3740 5102
rect 4172 5114 4200 5578
rect 4814 5468 5122 5477
rect 4814 5466 4820 5468
rect 4876 5466 4900 5468
rect 4956 5466 4980 5468
rect 5036 5466 5060 5468
rect 5116 5466 5122 5468
rect 4876 5414 4878 5466
rect 5058 5414 5060 5466
rect 4814 5412 4820 5414
rect 4876 5412 4900 5414
rect 4956 5412 4980 5414
rect 5036 5412 5060 5414
rect 5116 5412 5122 5414
rect 4814 5403 5122 5412
rect 4122 5086 4200 5114
rect 4066 5063 4122 5072
rect 3848 4924 4156 4933
rect 3848 4922 3854 4924
rect 3910 4922 3934 4924
rect 3990 4922 4014 4924
rect 4070 4922 4094 4924
rect 4150 4922 4156 4924
rect 3910 4870 3912 4922
rect 4092 4870 4094 4922
rect 3848 4868 3854 4870
rect 3910 4868 3934 4870
rect 3990 4868 4014 4870
rect 4070 4868 4094 4870
rect 4150 4868 4156 4870
rect 3848 4859 4156 4868
rect 3700 4616 3752 4622
rect 5184 4570 5212 6054
rect 5368 5302 5396 6598
rect 5828 6322 5856 6734
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6390 5948 6666
rect 6380 6390 6408 6938
rect 8312 6798 8340 7142
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5780 6012 6088 6021
rect 5780 6010 5786 6012
rect 5842 6010 5866 6012
rect 5922 6010 5946 6012
rect 6002 6010 6026 6012
rect 6082 6010 6088 6012
rect 5842 5958 5844 6010
rect 6024 5958 6026 6010
rect 5780 5956 5786 5958
rect 5842 5956 5866 5958
rect 5922 5956 5946 5958
rect 6002 5956 6026 5958
rect 6082 5956 6088 5958
rect 5780 5947 6088 5956
rect 6472 5642 6500 6598
rect 6746 6556 7054 6565
rect 6746 6554 6752 6556
rect 6808 6554 6832 6556
rect 6888 6554 6912 6556
rect 6968 6554 6992 6556
rect 7048 6554 7054 6556
rect 6808 6502 6810 6554
rect 6990 6502 6992 6554
rect 6746 6500 6752 6502
rect 6808 6500 6832 6502
rect 6888 6500 6912 6502
rect 6968 6500 6992 6502
rect 7048 6500 7054 6502
rect 6746 6491 7054 6500
rect 7116 6458 7144 6666
rect 8678 6556 8986 6565
rect 8678 6554 8684 6556
rect 8740 6554 8764 6556
rect 8820 6554 8844 6556
rect 8900 6554 8924 6556
rect 8980 6554 8986 6556
rect 8740 6502 8742 6554
rect 8922 6502 8924 6554
rect 8678 6500 8684 6502
rect 8740 6500 8764 6502
rect 8820 6500 8844 6502
rect 8900 6500 8924 6502
rect 8980 6500 8986 6502
rect 8678 6491 8986 6500
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6656 5574 6684 6258
rect 7116 5710 7144 6394
rect 7712 6012 8020 6021
rect 7712 6010 7718 6012
rect 7774 6010 7798 6012
rect 7854 6010 7878 6012
rect 7934 6010 7958 6012
rect 8014 6010 8020 6012
rect 7774 5958 7776 6010
rect 7956 5958 7958 6010
rect 7712 5956 7718 5958
rect 7774 5956 7798 5958
rect 7854 5956 7878 5958
rect 7934 5956 7958 5958
rect 8014 5956 8020 5958
rect 7712 5947 8020 5956
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 6746 5468 7054 5477
rect 6746 5466 6752 5468
rect 6808 5466 6832 5468
rect 6888 5466 6912 5468
rect 6968 5466 6992 5468
rect 7048 5466 7054 5468
rect 6808 5414 6810 5466
rect 6990 5414 6992 5466
rect 6746 5412 6752 5414
rect 6808 5412 6832 5414
rect 6888 5412 6912 5414
rect 6968 5412 6992 5414
rect 7048 5412 7054 5414
rect 6746 5403 7054 5412
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 3700 4558 3752 4564
rect 5092 4554 5212 4570
rect 5080 4548 5212 4554
rect 5132 4542 5212 4548
rect 5080 4490 5132 4496
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 1916 3836 2224 3845
rect 1916 3834 1922 3836
rect 1978 3834 2002 3836
rect 2058 3834 2082 3836
rect 2138 3834 2162 3836
rect 2218 3834 2224 3836
rect 1978 3782 1980 3834
rect 2160 3782 2162 3834
rect 1916 3780 1922 3782
rect 1978 3780 2002 3782
rect 2058 3780 2082 3782
rect 2138 3780 2162 3782
rect 2218 3780 2224 3782
rect 1916 3771 2224 3780
rect 1916 2748 2224 2757
rect 1916 2746 1922 2748
rect 1978 2746 2002 2748
rect 2058 2746 2082 2748
rect 2138 2746 2162 2748
rect 2218 2746 2224 2748
rect 1978 2694 1980 2746
rect 2160 2694 2162 2746
rect 1916 2692 1922 2694
rect 1978 2692 2002 2694
rect 2058 2692 2082 2694
rect 2138 2692 2162 2694
rect 2218 2692 2224 2694
rect 1916 2683 2224 2692
rect 2792 2446 2820 4422
rect 2882 4380 3190 4389
rect 2882 4378 2888 4380
rect 2944 4378 2968 4380
rect 3024 4378 3048 4380
rect 3104 4378 3128 4380
rect 3184 4378 3190 4380
rect 2944 4326 2946 4378
rect 3126 4326 3128 4378
rect 2882 4324 2888 4326
rect 2944 4324 2968 4326
rect 3024 4324 3048 4326
rect 3104 4324 3128 4326
rect 3184 4324 3190 4326
rect 2882 4315 3190 4324
rect 4814 4380 5122 4389
rect 4814 4378 4820 4380
rect 4876 4378 4900 4380
rect 4956 4378 4980 4380
rect 5036 4378 5060 4380
rect 5116 4378 5122 4380
rect 4876 4326 4878 4378
rect 5058 4326 5060 4378
rect 4814 4324 4820 4326
rect 4876 4324 4900 4326
rect 4956 4324 4980 4326
rect 5036 4324 5060 4326
rect 5116 4324 5122 4326
rect 4814 4315 5122 4324
rect 3848 3836 4156 3845
rect 3848 3834 3854 3836
rect 3910 3834 3934 3836
rect 3990 3834 4014 3836
rect 4070 3834 4094 3836
rect 4150 3834 4156 3836
rect 3910 3782 3912 3834
rect 4092 3782 4094 3834
rect 3848 3780 3854 3782
rect 3910 3780 3934 3782
rect 3990 3780 4014 3782
rect 4070 3780 4094 3782
rect 4150 3780 4156 3782
rect 3848 3771 4156 3780
rect 2882 3292 3190 3301
rect 2882 3290 2888 3292
rect 2944 3290 2968 3292
rect 3024 3290 3048 3292
rect 3104 3290 3128 3292
rect 3184 3290 3190 3292
rect 2944 3238 2946 3290
rect 3126 3238 3128 3290
rect 2882 3236 2888 3238
rect 2944 3236 2968 3238
rect 3024 3236 3048 3238
rect 3104 3236 3128 3238
rect 3184 3236 3190 3238
rect 2882 3227 3190 3236
rect 4814 3292 5122 3301
rect 4814 3290 4820 3292
rect 4876 3290 4900 3292
rect 4956 3290 4980 3292
rect 5036 3290 5060 3292
rect 5116 3290 5122 3292
rect 4876 3238 4878 3290
rect 5058 3238 5060 3290
rect 4814 3236 4820 3238
rect 4876 3236 4900 3238
rect 4956 3236 4980 3238
rect 5036 3236 5060 3238
rect 5116 3236 5122 3238
rect 4814 3227 5122 3236
rect 3848 2748 4156 2757
rect 3848 2746 3854 2748
rect 3910 2746 3934 2748
rect 3990 2746 4014 2748
rect 4070 2746 4094 2748
rect 4150 2746 4156 2748
rect 3910 2694 3912 2746
rect 4092 2694 4094 2746
rect 3848 2692 3854 2694
rect 3910 2692 3934 2694
rect 3990 2692 4014 2694
rect 4070 2692 4094 2694
rect 4150 2692 4156 2694
rect 3848 2683 4156 2692
rect 5368 2446 5396 4966
rect 5780 4924 6088 4933
rect 5780 4922 5786 4924
rect 5842 4922 5866 4924
rect 5922 4922 5946 4924
rect 6002 4922 6026 4924
rect 6082 4922 6088 4924
rect 5842 4870 5844 4922
rect 6024 4870 6026 4922
rect 5780 4868 5786 4870
rect 5842 4868 5866 4870
rect 5922 4868 5946 4870
rect 6002 4868 6026 4870
rect 6082 4868 6088 4870
rect 5780 4859 6088 4868
rect 7712 4924 8020 4933
rect 7712 4922 7718 4924
rect 7774 4922 7798 4924
rect 7854 4922 7878 4924
rect 7934 4922 7958 4924
rect 8014 4922 8020 4924
rect 7774 4870 7776 4922
rect 7956 4870 7958 4922
rect 7712 4868 7718 4870
rect 7774 4868 7798 4870
rect 7854 4868 7878 4870
rect 7934 4868 7958 4870
rect 8014 4868 8020 4870
rect 7712 4859 8020 4868
rect 6746 4380 7054 4389
rect 6746 4378 6752 4380
rect 6808 4378 6832 4380
rect 6888 4378 6912 4380
rect 6968 4378 6992 4380
rect 7048 4378 7054 4380
rect 6808 4326 6810 4378
rect 6990 4326 6992 4378
rect 6746 4324 6752 4326
rect 6808 4324 6832 4326
rect 6888 4324 6912 4326
rect 6968 4324 6992 4326
rect 7048 4324 7054 4326
rect 6746 4315 7054 4324
rect 5780 3836 6088 3845
rect 5780 3834 5786 3836
rect 5842 3834 5866 3836
rect 5922 3834 5946 3836
rect 6002 3834 6026 3836
rect 6082 3834 6088 3836
rect 5842 3782 5844 3834
rect 6024 3782 6026 3834
rect 5780 3780 5786 3782
rect 5842 3780 5866 3782
rect 5922 3780 5946 3782
rect 6002 3780 6026 3782
rect 6082 3780 6088 3782
rect 5780 3771 6088 3780
rect 7712 3836 8020 3845
rect 7712 3834 7718 3836
rect 7774 3834 7798 3836
rect 7854 3834 7878 3836
rect 7934 3834 7958 3836
rect 8014 3834 8020 3836
rect 7774 3782 7776 3834
rect 7956 3782 7958 3834
rect 7712 3780 7718 3782
rect 7774 3780 7798 3782
rect 7854 3780 7878 3782
rect 7934 3780 7958 3782
rect 8014 3780 8020 3782
rect 7712 3771 8020 3780
rect 6746 3292 7054 3301
rect 6746 3290 6752 3292
rect 6808 3290 6832 3292
rect 6888 3290 6912 3292
rect 6968 3290 6992 3292
rect 7048 3290 7054 3292
rect 6808 3238 6810 3290
rect 6990 3238 6992 3290
rect 6746 3236 6752 3238
rect 6808 3236 6832 3238
rect 6888 3236 6912 3238
rect 6968 3236 6992 3238
rect 7048 3236 7054 3238
rect 6746 3227 7054 3236
rect 5780 2748 6088 2757
rect 5780 2746 5786 2748
rect 5842 2746 5866 2748
rect 5922 2746 5946 2748
rect 6002 2746 6026 2748
rect 6082 2746 6088 2748
rect 5842 2694 5844 2746
rect 6024 2694 6026 2746
rect 5780 2692 5786 2694
rect 5842 2692 5866 2694
rect 5922 2692 5946 2694
rect 6002 2692 6026 2694
rect 6082 2692 6088 2694
rect 5780 2683 6088 2692
rect 7712 2748 8020 2757
rect 7712 2746 7718 2748
rect 7774 2746 7798 2748
rect 7854 2746 7878 2748
rect 7934 2746 7958 2748
rect 8014 2746 8020 2748
rect 7774 2694 7776 2746
rect 7956 2694 7958 2746
rect 7712 2692 7718 2694
rect 7774 2692 7798 2694
rect 7854 2692 7878 2694
rect 7934 2692 7958 2694
rect 8014 2692 8020 2694
rect 7712 2683 8020 2692
rect 8220 2446 8248 5510
rect 8678 5468 8986 5477
rect 8678 5466 8684 5468
rect 8740 5466 8764 5468
rect 8820 5466 8844 5468
rect 8900 5466 8924 5468
rect 8980 5466 8986 5468
rect 8740 5414 8742 5466
rect 8922 5414 8924 5466
rect 8678 5412 8684 5414
rect 8740 5412 8764 5414
rect 8820 5412 8844 5414
rect 8900 5412 8924 5414
rect 8980 5412 8986 5414
rect 8678 5403 8986 5412
rect 8678 4380 8986 4389
rect 8678 4378 8684 4380
rect 8740 4378 8764 4380
rect 8820 4378 8844 4380
rect 8900 4378 8924 4380
rect 8980 4378 8986 4380
rect 8740 4326 8742 4378
rect 8922 4326 8924 4378
rect 8678 4324 8684 4326
rect 8740 4324 8764 4326
rect 8820 4324 8844 4326
rect 8900 4324 8924 4326
rect 8980 4324 8986 4326
rect 8678 4315 8986 4324
rect 8678 3292 8986 3301
rect 8678 3290 8684 3292
rect 8740 3290 8764 3292
rect 8820 3290 8844 3292
rect 8900 3290 8924 3292
rect 8980 3290 8986 3292
rect 8740 3238 8742 3290
rect 8922 3238 8924 3290
rect 8678 3236 8684 3238
rect 8740 3236 8764 3238
rect 8820 3236 8844 3238
rect 8900 3236 8924 3238
rect 8980 3236 8986 3238
rect 8678 3227 8986 3236
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 1688 800 1716 2246
rect 2882 2204 3190 2213
rect 2882 2202 2888 2204
rect 2944 2202 2968 2204
rect 3024 2202 3048 2204
rect 3104 2202 3128 2204
rect 3184 2202 3190 2204
rect 2944 2150 2946 2202
rect 3126 2150 3128 2202
rect 2882 2148 2888 2150
rect 2944 2148 2968 2150
rect 3024 2148 3048 2150
rect 3104 2148 3128 2150
rect 3184 2148 3190 2150
rect 2882 2139 3190 2148
rect 4814 2204 5122 2213
rect 4814 2202 4820 2204
rect 4876 2202 4900 2204
rect 4956 2202 4980 2204
rect 5036 2202 5060 2204
rect 5116 2202 5122 2204
rect 4876 2150 4878 2202
rect 5058 2150 5060 2202
rect 4814 2148 4820 2150
rect 4876 2148 4900 2150
rect 4956 2148 4980 2150
rect 5036 2148 5060 2150
rect 5116 2148 5122 2150
rect 4814 2139 5122 2148
rect 5184 1170 5212 2246
rect 6746 2204 7054 2213
rect 6746 2202 6752 2204
rect 6808 2202 6832 2204
rect 6888 2202 6912 2204
rect 6968 2202 6992 2204
rect 7048 2202 7054 2204
rect 6808 2150 6810 2202
rect 6990 2150 6992 2202
rect 6746 2148 6752 2150
rect 6808 2148 6832 2150
rect 6888 2148 6912 2150
rect 6968 2148 6992 2150
rect 7048 2148 7054 2150
rect 6746 2139 7054 2148
rect 5000 1142 5212 1170
rect 5000 800 5028 1142
rect 8312 800 8340 2246
rect 8678 2204 8986 2213
rect 8678 2202 8684 2204
rect 8740 2202 8764 2204
rect 8820 2202 8844 2204
rect 8900 2202 8924 2204
rect 8980 2202 8986 2204
rect 8740 2150 8742 2202
rect 8922 2150 8924 2202
rect 8678 2148 8684 2150
rect 8740 2148 8764 2150
rect 8820 2148 8844 2150
rect 8900 2148 8924 2150
rect 8980 2148 8986 2150
rect 8678 2139 8986 2148
rect 1674 0 1730 800
rect 4986 0 5042 800
rect 8298 0 8354 800
<< via2 >>
rect 2888 7642 2944 7644
rect 2968 7642 3024 7644
rect 3048 7642 3104 7644
rect 3128 7642 3184 7644
rect 2888 7590 2934 7642
rect 2934 7590 2944 7642
rect 2968 7590 2998 7642
rect 2998 7590 3010 7642
rect 3010 7590 3024 7642
rect 3048 7590 3062 7642
rect 3062 7590 3074 7642
rect 3074 7590 3104 7642
rect 3128 7590 3138 7642
rect 3138 7590 3184 7642
rect 2888 7588 2944 7590
rect 2968 7588 3024 7590
rect 3048 7588 3104 7590
rect 3128 7588 3184 7590
rect 4820 7642 4876 7644
rect 4900 7642 4956 7644
rect 4980 7642 5036 7644
rect 5060 7642 5116 7644
rect 4820 7590 4866 7642
rect 4866 7590 4876 7642
rect 4900 7590 4930 7642
rect 4930 7590 4942 7642
rect 4942 7590 4956 7642
rect 4980 7590 4994 7642
rect 4994 7590 5006 7642
rect 5006 7590 5036 7642
rect 5060 7590 5070 7642
rect 5070 7590 5116 7642
rect 4820 7588 4876 7590
rect 4900 7588 4956 7590
rect 4980 7588 5036 7590
rect 5060 7588 5116 7590
rect 6752 7642 6808 7644
rect 6832 7642 6888 7644
rect 6912 7642 6968 7644
rect 6992 7642 7048 7644
rect 6752 7590 6798 7642
rect 6798 7590 6808 7642
rect 6832 7590 6862 7642
rect 6862 7590 6874 7642
rect 6874 7590 6888 7642
rect 6912 7590 6926 7642
rect 6926 7590 6938 7642
rect 6938 7590 6968 7642
rect 6992 7590 7002 7642
rect 7002 7590 7048 7642
rect 6752 7588 6808 7590
rect 6832 7588 6888 7590
rect 6912 7588 6968 7590
rect 6992 7588 7048 7590
rect 8684 7642 8740 7644
rect 8764 7642 8820 7644
rect 8844 7642 8900 7644
rect 8924 7642 8980 7644
rect 8684 7590 8730 7642
rect 8730 7590 8740 7642
rect 8764 7590 8794 7642
rect 8794 7590 8806 7642
rect 8806 7590 8820 7642
rect 8844 7590 8858 7642
rect 8858 7590 8870 7642
rect 8870 7590 8900 7642
rect 8924 7590 8934 7642
rect 8934 7590 8980 7642
rect 8684 7588 8740 7590
rect 8764 7588 8820 7590
rect 8844 7588 8900 7590
rect 8924 7588 8980 7590
rect 1922 7098 1978 7100
rect 2002 7098 2058 7100
rect 2082 7098 2138 7100
rect 2162 7098 2218 7100
rect 1922 7046 1968 7098
rect 1968 7046 1978 7098
rect 2002 7046 2032 7098
rect 2032 7046 2044 7098
rect 2044 7046 2058 7098
rect 2082 7046 2096 7098
rect 2096 7046 2108 7098
rect 2108 7046 2138 7098
rect 2162 7046 2172 7098
rect 2172 7046 2218 7098
rect 1922 7044 1978 7046
rect 2002 7044 2058 7046
rect 2082 7044 2138 7046
rect 2162 7044 2218 7046
rect 3854 7098 3910 7100
rect 3934 7098 3990 7100
rect 4014 7098 4070 7100
rect 4094 7098 4150 7100
rect 3854 7046 3900 7098
rect 3900 7046 3910 7098
rect 3934 7046 3964 7098
rect 3964 7046 3976 7098
rect 3976 7046 3990 7098
rect 4014 7046 4028 7098
rect 4028 7046 4040 7098
rect 4040 7046 4070 7098
rect 4094 7046 4104 7098
rect 4104 7046 4150 7098
rect 3854 7044 3910 7046
rect 3934 7044 3990 7046
rect 4014 7044 4070 7046
rect 4094 7044 4150 7046
rect 5786 7098 5842 7100
rect 5866 7098 5922 7100
rect 5946 7098 6002 7100
rect 6026 7098 6082 7100
rect 5786 7046 5832 7098
rect 5832 7046 5842 7098
rect 5866 7046 5896 7098
rect 5896 7046 5908 7098
rect 5908 7046 5922 7098
rect 5946 7046 5960 7098
rect 5960 7046 5972 7098
rect 5972 7046 6002 7098
rect 6026 7046 6036 7098
rect 6036 7046 6082 7098
rect 5786 7044 5842 7046
rect 5866 7044 5922 7046
rect 5946 7044 6002 7046
rect 6026 7044 6082 7046
rect 7718 7098 7774 7100
rect 7798 7098 7854 7100
rect 7878 7098 7934 7100
rect 7958 7098 8014 7100
rect 7718 7046 7764 7098
rect 7764 7046 7774 7098
rect 7798 7046 7828 7098
rect 7828 7046 7840 7098
rect 7840 7046 7854 7098
rect 7878 7046 7892 7098
rect 7892 7046 7904 7098
rect 7904 7046 7934 7098
rect 7958 7046 7968 7098
rect 7968 7046 8014 7098
rect 7718 7044 7774 7046
rect 7798 7044 7854 7046
rect 7878 7044 7934 7046
rect 7958 7044 8014 7046
rect 2888 6554 2944 6556
rect 2968 6554 3024 6556
rect 3048 6554 3104 6556
rect 3128 6554 3184 6556
rect 2888 6502 2934 6554
rect 2934 6502 2944 6554
rect 2968 6502 2998 6554
rect 2998 6502 3010 6554
rect 3010 6502 3024 6554
rect 3048 6502 3062 6554
rect 3062 6502 3074 6554
rect 3074 6502 3104 6554
rect 3128 6502 3138 6554
rect 3138 6502 3184 6554
rect 2888 6500 2944 6502
rect 2968 6500 3024 6502
rect 3048 6500 3104 6502
rect 3128 6500 3184 6502
rect 4820 6554 4876 6556
rect 4900 6554 4956 6556
rect 4980 6554 5036 6556
rect 5060 6554 5116 6556
rect 4820 6502 4866 6554
rect 4866 6502 4876 6554
rect 4900 6502 4930 6554
rect 4930 6502 4942 6554
rect 4942 6502 4956 6554
rect 4980 6502 4994 6554
rect 4994 6502 5006 6554
rect 5006 6502 5036 6554
rect 5060 6502 5070 6554
rect 5070 6502 5116 6554
rect 4820 6500 4876 6502
rect 4900 6500 4956 6502
rect 4980 6500 5036 6502
rect 5060 6500 5116 6502
rect 1922 6010 1978 6012
rect 2002 6010 2058 6012
rect 2082 6010 2138 6012
rect 2162 6010 2218 6012
rect 1922 5958 1968 6010
rect 1968 5958 1978 6010
rect 2002 5958 2032 6010
rect 2032 5958 2044 6010
rect 2044 5958 2058 6010
rect 2082 5958 2096 6010
rect 2096 5958 2108 6010
rect 2108 5958 2138 6010
rect 2162 5958 2172 6010
rect 2172 5958 2218 6010
rect 1922 5956 1978 5958
rect 2002 5956 2058 5958
rect 2082 5956 2138 5958
rect 2162 5956 2218 5958
rect 3854 6010 3910 6012
rect 3934 6010 3990 6012
rect 4014 6010 4070 6012
rect 4094 6010 4150 6012
rect 3854 5958 3900 6010
rect 3900 5958 3910 6010
rect 3934 5958 3964 6010
rect 3964 5958 3976 6010
rect 3976 5958 3990 6010
rect 4014 5958 4028 6010
rect 4028 5958 4040 6010
rect 4040 5958 4070 6010
rect 4094 5958 4104 6010
rect 4104 5958 4150 6010
rect 3854 5956 3910 5958
rect 3934 5956 3990 5958
rect 4014 5956 4070 5958
rect 4094 5956 4150 5958
rect 2888 5466 2944 5468
rect 2968 5466 3024 5468
rect 3048 5466 3104 5468
rect 3128 5466 3184 5468
rect 2888 5414 2934 5466
rect 2934 5414 2944 5466
rect 2968 5414 2998 5466
rect 2998 5414 3010 5466
rect 3010 5414 3024 5466
rect 3048 5414 3062 5466
rect 3062 5414 3074 5466
rect 3074 5414 3104 5466
rect 3128 5414 3138 5466
rect 3138 5414 3184 5466
rect 2888 5412 2944 5414
rect 2968 5412 3024 5414
rect 3048 5412 3104 5414
rect 3128 5412 3184 5414
rect 1922 4922 1978 4924
rect 2002 4922 2058 4924
rect 2082 4922 2138 4924
rect 2162 4922 2218 4924
rect 1922 4870 1968 4922
rect 1968 4870 1978 4922
rect 2002 4870 2032 4922
rect 2032 4870 2044 4922
rect 2044 4870 2058 4922
rect 2082 4870 2096 4922
rect 2096 4870 2108 4922
rect 2108 4870 2138 4922
rect 2162 4870 2172 4922
rect 2172 4870 2218 4922
rect 1922 4868 1978 4870
rect 2002 4868 2058 4870
rect 2082 4868 2138 4870
rect 2162 4868 2218 4870
rect 4066 5072 4122 5128
rect 4820 5466 4876 5468
rect 4900 5466 4956 5468
rect 4980 5466 5036 5468
rect 5060 5466 5116 5468
rect 4820 5414 4866 5466
rect 4866 5414 4876 5466
rect 4900 5414 4930 5466
rect 4930 5414 4942 5466
rect 4942 5414 4956 5466
rect 4980 5414 4994 5466
rect 4994 5414 5006 5466
rect 5006 5414 5036 5466
rect 5060 5414 5070 5466
rect 5070 5414 5116 5466
rect 4820 5412 4876 5414
rect 4900 5412 4956 5414
rect 4980 5412 5036 5414
rect 5060 5412 5116 5414
rect 3854 4922 3910 4924
rect 3934 4922 3990 4924
rect 4014 4922 4070 4924
rect 4094 4922 4150 4924
rect 3854 4870 3900 4922
rect 3900 4870 3910 4922
rect 3934 4870 3964 4922
rect 3964 4870 3976 4922
rect 3976 4870 3990 4922
rect 4014 4870 4028 4922
rect 4028 4870 4040 4922
rect 4040 4870 4070 4922
rect 4094 4870 4104 4922
rect 4104 4870 4150 4922
rect 3854 4868 3910 4870
rect 3934 4868 3990 4870
rect 4014 4868 4070 4870
rect 4094 4868 4150 4870
rect 5786 6010 5842 6012
rect 5866 6010 5922 6012
rect 5946 6010 6002 6012
rect 6026 6010 6082 6012
rect 5786 5958 5832 6010
rect 5832 5958 5842 6010
rect 5866 5958 5896 6010
rect 5896 5958 5908 6010
rect 5908 5958 5922 6010
rect 5946 5958 5960 6010
rect 5960 5958 5972 6010
rect 5972 5958 6002 6010
rect 6026 5958 6036 6010
rect 6036 5958 6082 6010
rect 5786 5956 5842 5958
rect 5866 5956 5922 5958
rect 5946 5956 6002 5958
rect 6026 5956 6082 5958
rect 6752 6554 6808 6556
rect 6832 6554 6888 6556
rect 6912 6554 6968 6556
rect 6992 6554 7048 6556
rect 6752 6502 6798 6554
rect 6798 6502 6808 6554
rect 6832 6502 6862 6554
rect 6862 6502 6874 6554
rect 6874 6502 6888 6554
rect 6912 6502 6926 6554
rect 6926 6502 6938 6554
rect 6938 6502 6968 6554
rect 6992 6502 7002 6554
rect 7002 6502 7048 6554
rect 6752 6500 6808 6502
rect 6832 6500 6888 6502
rect 6912 6500 6968 6502
rect 6992 6500 7048 6502
rect 8684 6554 8740 6556
rect 8764 6554 8820 6556
rect 8844 6554 8900 6556
rect 8924 6554 8980 6556
rect 8684 6502 8730 6554
rect 8730 6502 8740 6554
rect 8764 6502 8794 6554
rect 8794 6502 8806 6554
rect 8806 6502 8820 6554
rect 8844 6502 8858 6554
rect 8858 6502 8870 6554
rect 8870 6502 8900 6554
rect 8924 6502 8934 6554
rect 8934 6502 8980 6554
rect 8684 6500 8740 6502
rect 8764 6500 8820 6502
rect 8844 6500 8900 6502
rect 8924 6500 8980 6502
rect 7718 6010 7774 6012
rect 7798 6010 7854 6012
rect 7878 6010 7934 6012
rect 7958 6010 8014 6012
rect 7718 5958 7764 6010
rect 7764 5958 7774 6010
rect 7798 5958 7828 6010
rect 7828 5958 7840 6010
rect 7840 5958 7854 6010
rect 7878 5958 7892 6010
rect 7892 5958 7904 6010
rect 7904 5958 7934 6010
rect 7958 5958 7968 6010
rect 7968 5958 8014 6010
rect 7718 5956 7774 5958
rect 7798 5956 7854 5958
rect 7878 5956 7934 5958
rect 7958 5956 8014 5958
rect 6752 5466 6808 5468
rect 6832 5466 6888 5468
rect 6912 5466 6968 5468
rect 6992 5466 7048 5468
rect 6752 5414 6798 5466
rect 6798 5414 6808 5466
rect 6832 5414 6862 5466
rect 6862 5414 6874 5466
rect 6874 5414 6888 5466
rect 6912 5414 6926 5466
rect 6926 5414 6938 5466
rect 6938 5414 6968 5466
rect 6992 5414 7002 5466
rect 7002 5414 7048 5466
rect 6752 5412 6808 5414
rect 6832 5412 6888 5414
rect 6912 5412 6968 5414
rect 6992 5412 7048 5414
rect 1922 3834 1978 3836
rect 2002 3834 2058 3836
rect 2082 3834 2138 3836
rect 2162 3834 2218 3836
rect 1922 3782 1968 3834
rect 1968 3782 1978 3834
rect 2002 3782 2032 3834
rect 2032 3782 2044 3834
rect 2044 3782 2058 3834
rect 2082 3782 2096 3834
rect 2096 3782 2108 3834
rect 2108 3782 2138 3834
rect 2162 3782 2172 3834
rect 2172 3782 2218 3834
rect 1922 3780 1978 3782
rect 2002 3780 2058 3782
rect 2082 3780 2138 3782
rect 2162 3780 2218 3782
rect 1922 2746 1978 2748
rect 2002 2746 2058 2748
rect 2082 2746 2138 2748
rect 2162 2746 2218 2748
rect 1922 2694 1968 2746
rect 1968 2694 1978 2746
rect 2002 2694 2032 2746
rect 2032 2694 2044 2746
rect 2044 2694 2058 2746
rect 2082 2694 2096 2746
rect 2096 2694 2108 2746
rect 2108 2694 2138 2746
rect 2162 2694 2172 2746
rect 2172 2694 2218 2746
rect 1922 2692 1978 2694
rect 2002 2692 2058 2694
rect 2082 2692 2138 2694
rect 2162 2692 2218 2694
rect 2888 4378 2944 4380
rect 2968 4378 3024 4380
rect 3048 4378 3104 4380
rect 3128 4378 3184 4380
rect 2888 4326 2934 4378
rect 2934 4326 2944 4378
rect 2968 4326 2998 4378
rect 2998 4326 3010 4378
rect 3010 4326 3024 4378
rect 3048 4326 3062 4378
rect 3062 4326 3074 4378
rect 3074 4326 3104 4378
rect 3128 4326 3138 4378
rect 3138 4326 3184 4378
rect 2888 4324 2944 4326
rect 2968 4324 3024 4326
rect 3048 4324 3104 4326
rect 3128 4324 3184 4326
rect 4820 4378 4876 4380
rect 4900 4378 4956 4380
rect 4980 4378 5036 4380
rect 5060 4378 5116 4380
rect 4820 4326 4866 4378
rect 4866 4326 4876 4378
rect 4900 4326 4930 4378
rect 4930 4326 4942 4378
rect 4942 4326 4956 4378
rect 4980 4326 4994 4378
rect 4994 4326 5006 4378
rect 5006 4326 5036 4378
rect 5060 4326 5070 4378
rect 5070 4326 5116 4378
rect 4820 4324 4876 4326
rect 4900 4324 4956 4326
rect 4980 4324 5036 4326
rect 5060 4324 5116 4326
rect 3854 3834 3910 3836
rect 3934 3834 3990 3836
rect 4014 3834 4070 3836
rect 4094 3834 4150 3836
rect 3854 3782 3900 3834
rect 3900 3782 3910 3834
rect 3934 3782 3964 3834
rect 3964 3782 3976 3834
rect 3976 3782 3990 3834
rect 4014 3782 4028 3834
rect 4028 3782 4040 3834
rect 4040 3782 4070 3834
rect 4094 3782 4104 3834
rect 4104 3782 4150 3834
rect 3854 3780 3910 3782
rect 3934 3780 3990 3782
rect 4014 3780 4070 3782
rect 4094 3780 4150 3782
rect 2888 3290 2944 3292
rect 2968 3290 3024 3292
rect 3048 3290 3104 3292
rect 3128 3290 3184 3292
rect 2888 3238 2934 3290
rect 2934 3238 2944 3290
rect 2968 3238 2998 3290
rect 2998 3238 3010 3290
rect 3010 3238 3024 3290
rect 3048 3238 3062 3290
rect 3062 3238 3074 3290
rect 3074 3238 3104 3290
rect 3128 3238 3138 3290
rect 3138 3238 3184 3290
rect 2888 3236 2944 3238
rect 2968 3236 3024 3238
rect 3048 3236 3104 3238
rect 3128 3236 3184 3238
rect 4820 3290 4876 3292
rect 4900 3290 4956 3292
rect 4980 3290 5036 3292
rect 5060 3290 5116 3292
rect 4820 3238 4866 3290
rect 4866 3238 4876 3290
rect 4900 3238 4930 3290
rect 4930 3238 4942 3290
rect 4942 3238 4956 3290
rect 4980 3238 4994 3290
rect 4994 3238 5006 3290
rect 5006 3238 5036 3290
rect 5060 3238 5070 3290
rect 5070 3238 5116 3290
rect 4820 3236 4876 3238
rect 4900 3236 4956 3238
rect 4980 3236 5036 3238
rect 5060 3236 5116 3238
rect 3854 2746 3910 2748
rect 3934 2746 3990 2748
rect 4014 2746 4070 2748
rect 4094 2746 4150 2748
rect 3854 2694 3900 2746
rect 3900 2694 3910 2746
rect 3934 2694 3964 2746
rect 3964 2694 3976 2746
rect 3976 2694 3990 2746
rect 4014 2694 4028 2746
rect 4028 2694 4040 2746
rect 4040 2694 4070 2746
rect 4094 2694 4104 2746
rect 4104 2694 4150 2746
rect 3854 2692 3910 2694
rect 3934 2692 3990 2694
rect 4014 2692 4070 2694
rect 4094 2692 4150 2694
rect 5786 4922 5842 4924
rect 5866 4922 5922 4924
rect 5946 4922 6002 4924
rect 6026 4922 6082 4924
rect 5786 4870 5832 4922
rect 5832 4870 5842 4922
rect 5866 4870 5896 4922
rect 5896 4870 5908 4922
rect 5908 4870 5922 4922
rect 5946 4870 5960 4922
rect 5960 4870 5972 4922
rect 5972 4870 6002 4922
rect 6026 4870 6036 4922
rect 6036 4870 6082 4922
rect 5786 4868 5842 4870
rect 5866 4868 5922 4870
rect 5946 4868 6002 4870
rect 6026 4868 6082 4870
rect 7718 4922 7774 4924
rect 7798 4922 7854 4924
rect 7878 4922 7934 4924
rect 7958 4922 8014 4924
rect 7718 4870 7764 4922
rect 7764 4870 7774 4922
rect 7798 4870 7828 4922
rect 7828 4870 7840 4922
rect 7840 4870 7854 4922
rect 7878 4870 7892 4922
rect 7892 4870 7904 4922
rect 7904 4870 7934 4922
rect 7958 4870 7968 4922
rect 7968 4870 8014 4922
rect 7718 4868 7774 4870
rect 7798 4868 7854 4870
rect 7878 4868 7934 4870
rect 7958 4868 8014 4870
rect 6752 4378 6808 4380
rect 6832 4378 6888 4380
rect 6912 4378 6968 4380
rect 6992 4378 7048 4380
rect 6752 4326 6798 4378
rect 6798 4326 6808 4378
rect 6832 4326 6862 4378
rect 6862 4326 6874 4378
rect 6874 4326 6888 4378
rect 6912 4326 6926 4378
rect 6926 4326 6938 4378
rect 6938 4326 6968 4378
rect 6992 4326 7002 4378
rect 7002 4326 7048 4378
rect 6752 4324 6808 4326
rect 6832 4324 6888 4326
rect 6912 4324 6968 4326
rect 6992 4324 7048 4326
rect 5786 3834 5842 3836
rect 5866 3834 5922 3836
rect 5946 3834 6002 3836
rect 6026 3834 6082 3836
rect 5786 3782 5832 3834
rect 5832 3782 5842 3834
rect 5866 3782 5896 3834
rect 5896 3782 5908 3834
rect 5908 3782 5922 3834
rect 5946 3782 5960 3834
rect 5960 3782 5972 3834
rect 5972 3782 6002 3834
rect 6026 3782 6036 3834
rect 6036 3782 6082 3834
rect 5786 3780 5842 3782
rect 5866 3780 5922 3782
rect 5946 3780 6002 3782
rect 6026 3780 6082 3782
rect 7718 3834 7774 3836
rect 7798 3834 7854 3836
rect 7878 3834 7934 3836
rect 7958 3834 8014 3836
rect 7718 3782 7764 3834
rect 7764 3782 7774 3834
rect 7798 3782 7828 3834
rect 7828 3782 7840 3834
rect 7840 3782 7854 3834
rect 7878 3782 7892 3834
rect 7892 3782 7904 3834
rect 7904 3782 7934 3834
rect 7958 3782 7968 3834
rect 7968 3782 8014 3834
rect 7718 3780 7774 3782
rect 7798 3780 7854 3782
rect 7878 3780 7934 3782
rect 7958 3780 8014 3782
rect 6752 3290 6808 3292
rect 6832 3290 6888 3292
rect 6912 3290 6968 3292
rect 6992 3290 7048 3292
rect 6752 3238 6798 3290
rect 6798 3238 6808 3290
rect 6832 3238 6862 3290
rect 6862 3238 6874 3290
rect 6874 3238 6888 3290
rect 6912 3238 6926 3290
rect 6926 3238 6938 3290
rect 6938 3238 6968 3290
rect 6992 3238 7002 3290
rect 7002 3238 7048 3290
rect 6752 3236 6808 3238
rect 6832 3236 6888 3238
rect 6912 3236 6968 3238
rect 6992 3236 7048 3238
rect 5786 2746 5842 2748
rect 5866 2746 5922 2748
rect 5946 2746 6002 2748
rect 6026 2746 6082 2748
rect 5786 2694 5832 2746
rect 5832 2694 5842 2746
rect 5866 2694 5896 2746
rect 5896 2694 5908 2746
rect 5908 2694 5922 2746
rect 5946 2694 5960 2746
rect 5960 2694 5972 2746
rect 5972 2694 6002 2746
rect 6026 2694 6036 2746
rect 6036 2694 6082 2746
rect 5786 2692 5842 2694
rect 5866 2692 5922 2694
rect 5946 2692 6002 2694
rect 6026 2692 6082 2694
rect 7718 2746 7774 2748
rect 7798 2746 7854 2748
rect 7878 2746 7934 2748
rect 7958 2746 8014 2748
rect 7718 2694 7764 2746
rect 7764 2694 7774 2746
rect 7798 2694 7828 2746
rect 7828 2694 7840 2746
rect 7840 2694 7854 2746
rect 7878 2694 7892 2746
rect 7892 2694 7904 2746
rect 7904 2694 7934 2746
rect 7958 2694 7968 2746
rect 7968 2694 8014 2746
rect 7718 2692 7774 2694
rect 7798 2692 7854 2694
rect 7878 2692 7934 2694
rect 7958 2692 8014 2694
rect 8684 5466 8740 5468
rect 8764 5466 8820 5468
rect 8844 5466 8900 5468
rect 8924 5466 8980 5468
rect 8684 5414 8730 5466
rect 8730 5414 8740 5466
rect 8764 5414 8794 5466
rect 8794 5414 8806 5466
rect 8806 5414 8820 5466
rect 8844 5414 8858 5466
rect 8858 5414 8870 5466
rect 8870 5414 8900 5466
rect 8924 5414 8934 5466
rect 8934 5414 8980 5466
rect 8684 5412 8740 5414
rect 8764 5412 8820 5414
rect 8844 5412 8900 5414
rect 8924 5412 8980 5414
rect 8684 4378 8740 4380
rect 8764 4378 8820 4380
rect 8844 4378 8900 4380
rect 8924 4378 8980 4380
rect 8684 4326 8730 4378
rect 8730 4326 8740 4378
rect 8764 4326 8794 4378
rect 8794 4326 8806 4378
rect 8806 4326 8820 4378
rect 8844 4326 8858 4378
rect 8858 4326 8870 4378
rect 8870 4326 8900 4378
rect 8924 4326 8934 4378
rect 8934 4326 8980 4378
rect 8684 4324 8740 4326
rect 8764 4324 8820 4326
rect 8844 4324 8900 4326
rect 8924 4324 8980 4326
rect 8684 3290 8740 3292
rect 8764 3290 8820 3292
rect 8844 3290 8900 3292
rect 8924 3290 8980 3292
rect 8684 3238 8730 3290
rect 8730 3238 8740 3290
rect 8764 3238 8794 3290
rect 8794 3238 8806 3290
rect 8806 3238 8820 3290
rect 8844 3238 8858 3290
rect 8858 3238 8870 3290
rect 8870 3238 8900 3290
rect 8924 3238 8934 3290
rect 8934 3238 8980 3290
rect 8684 3236 8740 3238
rect 8764 3236 8820 3238
rect 8844 3236 8900 3238
rect 8924 3236 8980 3238
rect 2888 2202 2944 2204
rect 2968 2202 3024 2204
rect 3048 2202 3104 2204
rect 3128 2202 3184 2204
rect 2888 2150 2934 2202
rect 2934 2150 2944 2202
rect 2968 2150 2998 2202
rect 2998 2150 3010 2202
rect 3010 2150 3024 2202
rect 3048 2150 3062 2202
rect 3062 2150 3074 2202
rect 3074 2150 3104 2202
rect 3128 2150 3138 2202
rect 3138 2150 3184 2202
rect 2888 2148 2944 2150
rect 2968 2148 3024 2150
rect 3048 2148 3104 2150
rect 3128 2148 3184 2150
rect 4820 2202 4876 2204
rect 4900 2202 4956 2204
rect 4980 2202 5036 2204
rect 5060 2202 5116 2204
rect 4820 2150 4866 2202
rect 4866 2150 4876 2202
rect 4900 2150 4930 2202
rect 4930 2150 4942 2202
rect 4942 2150 4956 2202
rect 4980 2150 4994 2202
rect 4994 2150 5006 2202
rect 5006 2150 5036 2202
rect 5060 2150 5070 2202
rect 5070 2150 5116 2202
rect 4820 2148 4876 2150
rect 4900 2148 4956 2150
rect 4980 2148 5036 2150
rect 5060 2148 5116 2150
rect 6752 2202 6808 2204
rect 6832 2202 6888 2204
rect 6912 2202 6968 2204
rect 6992 2202 7048 2204
rect 6752 2150 6798 2202
rect 6798 2150 6808 2202
rect 6832 2150 6862 2202
rect 6862 2150 6874 2202
rect 6874 2150 6888 2202
rect 6912 2150 6926 2202
rect 6926 2150 6938 2202
rect 6938 2150 6968 2202
rect 6992 2150 7002 2202
rect 7002 2150 7048 2202
rect 6752 2148 6808 2150
rect 6832 2148 6888 2150
rect 6912 2148 6968 2150
rect 6992 2148 7048 2150
rect 8684 2202 8740 2204
rect 8764 2202 8820 2204
rect 8844 2202 8900 2204
rect 8924 2202 8980 2204
rect 8684 2150 8730 2202
rect 8730 2150 8740 2202
rect 8764 2150 8794 2202
rect 8794 2150 8806 2202
rect 8806 2150 8820 2202
rect 8844 2150 8858 2202
rect 8858 2150 8870 2202
rect 8870 2150 8900 2202
rect 8924 2150 8934 2202
rect 8934 2150 8980 2202
rect 8684 2148 8740 2150
rect 8764 2148 8820 2150
rect 8844 2148 8900 2150
rect 8924 2148 8980 2150
<< metal3 >>
rect 2878 7648 3194 7649
rect 2878 7584 2884 7648
rect 2948 7584 2964 7648
rect 3028 7584 3044 7648
rect 3108 7584 3124 7648
rect 3188 7584 3194 7648
rect 2878 7583 3194 7584
rect 4810 7648 5126 7649
rect 4810 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5126 7648
rect 4810 7583 5126 7584
rect 6742 7648 7058 7649
rect 6742 7584 6748 7648
rect 6812 7584 6828 7648
rect 6892 7584 6908 7648
rect 6972 7584 6988 7648
rect 7052 7584 7058 7648
rect 6742 7583 7058 7584
rect 8674 7648 8990 7649
rect 8674 7584 8680 7648
rect 8744 7584 8760 7648
rect 8824 7584 8840 7648
rect 8904 7584 8920 7648
rect 8984 7584 8990 7648
rect 8674 7583 8990 7584
rect 1912 7104 2228 7105
rect 1912 7040 1918 7104
rect 1982 7040 1998 7104
rect 2062 7040 2078 7104
rect 2142 7040 2158 7104
rect 2222 7040 2228 7104
rect 1912 7039 2228 7040
rect 3844 7104 4160 7105
rect 3844 7040 3850 7104
rect 3914 7040 3930 7104
rect 3994 7040 4010 7104
rect 4074 7040 4090 7104
rect 4154 7040 4160 7104
rect 3844 7039 4160 7040
rect 5776 7104 6092 7105
rect 5776 7040 5782 7104
rect 5846 7040 5862 7104
rect 5926 7040 5942 7104
rect 6006 7040 6022 7104
rect 6086 7040 6092 7104
rect 5776 7039 6092 7040
rect 7708 7104 8024 7105
rect 7708 7040 7714 7104
rect 7778 7040 7794 7104
rect 7858 7040 7874 7104
rect 7938 7040 7954 7104
rect 8018 7040 8024 7104
rect 7708 7039 8024 7040
rect 2878 6560 3194 6561
rect 2878 6496 2884 6560
rect 2948 6496 2964 6560
rect 3028 6496 3044 6560
rect 3108 6496 3124 6560
rect 3188 6496 3194 6560
rect 2878 6495 3194 6496
rect 4810 6560 5126 6561
rect 4810 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5126 6560
rect 4810 6495 5126 6496
rect 6742 6560 7058 6561
rect 6742 6496 6748 6560
rect 6812 6496 6828 6560
rect 6892 6496 6908 6560
rect 6972 6496 6988 6560
rect 7052 6496 7058 6560
rect 6742 6495 7058 6496
rect 8674 6560 8990 6561
rect 8674 6496 8680 6560
rect 8744 6496 8760 6560
rect 8824 6496 8840 6560
rect 8904 6496 8920 6560
rect 8984 6496 8990 6560
rect 8674 6495 8990 6496
rect 1912 6016 2228 6017
rect 1912 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2228 6016
rect 1912 5951 2228 5952
rect 3844 6016 4160 6017
rect 3844 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4160 6016
rect 3844 5951 4160 5952
rect 5776 6016 6092 6017
rect 5776 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6092 6016
rect 5776 5951 6092 5952
rect 7708 6016 8024 6017
rect 7708 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8024 6016
rect 7708 5951 8024 5952
rect 2878 5472 3194 5473
rect 2878 5408 2884 5472
rect 2948 5408 2964 5472
rect 3028 5408 3044 5472
rect 3108 5408 3124 5472
rect 3188 5408 3194 5472
rect 2878 5407 3194 5408
rect 4810 5472 5126 5473
rect 4810 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5126 5472
rect 4810 5407 5126 5408
rect 6742 5472 7058 5473
rect 6742 5408 6748 5472
rect 6812 5408 6828 5472
rect 6892 5408 6908 5472
rect 6972 5408 6988 5472
rect 7052 5408 7058 5472
rect 6742 5407 7058 5408
rect 8674 5472 8990 5473
rect 8674 5408 8680 5472
rect 8744 5408 8760 5472
rect 8824 5408 8840 5472
rect 8904 5408 8920 5472
rect 8984 5408 8990 5472
rect 8674 5407 8990 5408
rect 4061 5130 4127 5133
rect 1718 5128 4127 5130
rect 1718 5072 4066 5128
rect 4122 5072 4127 5128
rect 1718 5070 4127 5072
rect 0 4994 800 5024
rect 1718 4994 1778 5070
rect 4061 5067 4127 5070
rect 0 4934 1778 4994
rect 0 4904 800 4934
rect 1912 4928 2228 4929
rect 1912 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2228 4928
rect 1912 4863 2228 4864
rect 3844 4928 4160 4929
rect 3844 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4160 4928
rect 3844 4863 4160 4864
rect 5776 4928 6092 4929
rect 5776 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6092 4928
rect 5776 4863 6092 4864
rect 7708 4928 8024 4929
rect 7708 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8024 4928
rect 7708 4863 8024 4864
rect 2878 4384 3194 4385
rect 2878 4320 2884 4384
rect 2948 4320 2964 4384
rect 3028 4320 3044 4384
rect 3108 4320 3124 4384
rect 3188 4320 3194 4384
rect 2878 4319 3194 4320
rect 4810 4384 5126 4385
rect 4810 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5126 4384
rect 4810 4319 5126 4320
rect 6742 4384 7058 4385
rect 6742 4320 6748 4384
rect 6812 4320 6828 4384
rect 6892 4320 6908 4384
rect 6972 4320 6988 4384
rect 7052 4320 7058 4384
rect 6742 4319 7058 4320
rect 8674 4384 8990 4385
rect 8674 4320 8680 4384
rect 8744 4320 8760 4384
rect 8824 4320 8840 4384
rect 8904 4320 8920 4384
rect 8984 4320 8990 4384
rect 8674 4319 8990 4320
rect 1912 3840 2228 3841
rect 1912 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2228 3840
rect 1912 3775 2228 3776
rect 3844 3840 4160 3841
rect 3844 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4160 3840
rect 3844 3775 4160 3776
rect 5776 3840 6092 3841
rect 5776 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6092 3840
rect 5776 3775 6092 3776
rect 7708 3840 8024 3841
rect 7708 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8024 3840
rect 7708 3775 8024 3776
rect 2878 3296 3194 3297
rect 2878 3232 2884 3296
rect 2948 3232 2964 3296
rect 3028 3232 3044 3296
rect 3108 3232 3124 3296
rect 3188 3232 3194 3296
rect 2878 3231 3194 3232
rect 4810 3296 5126 3297
rect 4810 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5126 3296
rect 4810 3231 5126 3232
rect 6742 3296 7058 3297
rect 6742 3232 6748 3296
rect 6812 3232 6828 3296
rect 6892 3232 6908 3296
rect 6972 3232 6988 3296
rect 7052 3232 7058 3296
rect 6742 3231 7058 3232
rect 8674 3296 8990 3297
rect 8674 3232 8680 3296
rect 8744 3232 8760 3296
rect 8824 3232 8840 3296
rect 8904 3232 8920 3296
rect 8984 3232 8990 3296
rect 8674 3231 8990 3232
rect 1912 2752 2228 2753
rect 1912 2688 1918 2752
rect 1982 2688 1998 2752
rect 2062 2688 2078 2752
rect 2142 2688 2158 2752
rect 2222 2688 2228 2752
rect 1912 2687 2228 2688
rect 3844 2752 4160 2753
rect 3844 2688 3850 2752
rect 3914 2688 3930 2752
rect 3994 2688 4010 2752
rect 4074 2688 4090 2752
rect 4154 2688 4160 2752
rect 3844 2687 4160 2688
rect 5776 2752 6092 2753
rect 5776 2688 5782 2752
rect 5846 2688 5862 2752
rect 5926 2688 5942 2752
rect 6006 2688 6022 2752
rect 6086 2688 6092 2752
rect 5776 2687 6092 2688
rect 7708 2752 8024 2753
rect 7708 2688 7714 2752
rect 7778 2688 7794 2752
rect 7858 2688 7874 2752
rect 7938 2688 7954 2752
rect 8018 2688 8024 2752
rect 7708 2687 8024 2688
rect 2878 2208 3194 2209
rect 2878 2144 2884 2208
rect 2948 2144 2964 2208
rect 3028 2144 3044 2208
rect 3108 2144 3124 2208
rect 3188 2144 3194 2208
rect 2878 2143 3194 2144
rect 4810 2208 5126 2209
rect 4810 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5126 2208
rect 4810 2143 5126 2144
rect 6742 2208 7058 2209
rect 6742 2144 6748 2208
rect 6812 2144 6828 2208
rect 6892 2144 6908 2208
rect 6972 2144 6988 2208
rect 7052 2144 7058 2208
rect 6742 2143 7058 2144
rect 8674 2208 8990 2209
rect 8674 2144 8680 2208
rect 8744 2144 8760 2208
rect 8824 2144 8840 2208
rect 8904 2144 8920 2208
rect 8984 2144 8990 2208
rect 8674 2143 8990 2144
<< via3 >>
rect 2884 7644 2948 7648
rect 2884 7588 2888 7644
rect 2888 7588 2944 7644
rect 2944 7588 2948 7644
rect 2884 7584 2948 7588
rect 2964 7644 3028 7648
rect 2964 7588 2968 7644
rect 2968 7588 3024 7644
rect 3024 7588 3028 7644
rect 2964 7584 3028 7588
rect 3044 7644 3108 7648
rect 3044 7588 3048 7644
rect 3048 7588 3104 7644
rect 3104 7588 3108 7644
rect 3044 7584 3108 7588
rect 3124 7644 3188 7648
rect 3124 7588 3128 7644
rect 3128 7588 3184 7644
rect 3184 7588 3188 7644
rect 3124 7584 3188 7588
rect 4816 7644 4880 7648
rect 4816 7588 4820 7644
rect 4820 7588 4876 7644
rect 4876 7588 4880 7644
rect 4816 7584 4880 7588
rect 4896 7644 4960 7648
rect 4896 7588 4900 7644
rect 4900 7588 4956 7644
rect 4956 7588 4960 7644
rect 4896 7584 4960 7588
rect 4976 7644 5040 7648
rect 4976 7588 4980 7644
rect 4980 7588 5036 7644
rect 5036 7588 5040 7644
rect 4976 7584 5040 7588
rect 5056 7644 5120 7648
rect 5056 7588 5060 7644
rect 5060 7588 5116 7644
rect 5116 7588 5120 7644
rect 5056 7584 5120 7588
rect 6748 7644 6812 7648
rect 6748 7588 6752 7644
rect 6752 7588 6808 7644
rect 6808 7588 6812 7644
rect 6748 7584 6812 7588
rect 6828 7644 6892 7648
rect 6828 7588 6832 7644
rect 6832 7588 6888 7644
rect 6888 7588 6892 7644
rect 6828 7584 6892 7588
rect 6908 7644 6972 7648
rect 6908 7588 6912 7644
rect 6912 7588 6968 7644
rect 6968 7588 6972 7644
rect 6908 7584 6972 7588
rect 6988 7644 7052 7648
rect 6988 7588 6992 7644
rect 6992 7588 7048 7644
rect 7048 7588 7052 7644
rect 6988 7584 7052 7588
rect 8680 7644 8744 7648
rect 8680 7588 8684 7644
rect 8684 7588 8740 7644
rect 8740 7588 8744 7644
rect 8680 7584 8744 7588
rect 8760 7644 8824 7648
rect 8760 7588 8764 7644
rect 8764 7588 8820 7644
rect 8820 7588 8824 7644
rect 8760 7584 8824 7588
rect 8840 7644 8904 7648
rect 8840 7588 8844 7644
rect 8844 7588 8900 7644
rect 8900 7588 8904 7644
rect 8840 7584 8904 7588
rect 8920 7644 8984 7648
rect 8920 7588 8924 7644
rect 8924 7588 8980 7644
rect 8980 7588 8984 7644
rect 8920 7584 8984 7588
rect 1918 7100 1982 7104
rect 1918 7044 1922 7100
rect 1922 7044 1978 7100
rect 1978 7044 1982 7100
rect 1918 7040 1982 7044
rect 1998 7100 2062 7104
rect 1998 7044 2002 7100
rect 2002 7044 2058 7100
rect 2058 7044 2062 7100
rect 1998 7040 2062 7044
rect 2078 7100 2142 7104
rect 2078 7044 2082 7100
rect 2082 7044 2138 7100
rect 2138 7044 2142 7100
rect 2078 7040 2142 7044
rect 2158 7100 2222 7104
rect 2158 7044 2162 7100
rect 2162 7044 2218 7100
rect 2218 7044 2222 7100
rect 2158 7040 2222 7044
rect 3850 7100 3914 7104
rect 3850 7044 3854 7100
rect 3854 7044 3910 7100
rect 3910 7044 3914 7100
rect 3850 7040 3914 7044
rect 3930 7100 3994 7104
rect 3930 7044 3934 7100
rect 3934 7044 3990 7100
rect 3990 7044 3994 7100
rect 3930 7040 3994 7044
rect 4010 7100 4074 7104
rect 4010 7044 4014 7100
rect 4014 7044 4070 7100
rect 4070 7044 4074 7100
rect 4010 7040 4074 7044
rect 4090 7100 4154 7104
rect 4090 7044 4094 7100
rect 4094 7044 4150 7100
rect 4150 7044 4154 7100
rect 4090 7040 4154 7044
rect 5782 7100 5846 7104
rect 5782 7044 5786 7100
rect 5786 7044 5842 7100
rect 5842 7044 5846 7100
rect 5782 7040 5846 7044
rect 5862 7100 5926 7104
rect 5862 7044 5866 7100
rect 5866 7044 5922 7100
rect 5922 7044 5926 7100
rect 5862 7040 5926 7044
rect 5942 7100 6006 7104
rect 5942 7044 5946 7100
rect 5946 7044 6002 7100
rect 6002 7044 6006 7100
rect 5942 7040 6006 7044
rect 6022 7100 6086 7104
rect 6022 7044 6026 7100
rect 6026 7044 6082 7100
rect 6082 7044 6086 7100
rect 6022 7040 6086 7044
rect 7714 7100 7778 7104
rect 7714 7044 7718 7100
rect 7718 7044 7774 7100
rect 7774 7044 7778 7100
rect 7714 7040 7778 7044
rect 7794 7100 7858 7104
rect 7794 7044 7798 7100
rect 7798 7044 7854 7100
rect 7854 7044 7858 7100
rect 7794 7040 7858 7044
rect 7874 7100 7938 7104
rect 7874 7044 7878 7100
rect 7878 7044 7934 7100
rect 7934 7044 7938 7100
rect 7874 7040 7938 7044
rect 7954 7100 8018 7104
rect 7954 7044 7958 7100
rect 7958 7044 8014 7100
rect 8014 7044 8018 7100
rect 7954 7040 8018 7044
rect 2884 6556 2948 6560
rect 2884 6500 2888 6556
rect 2888 6500 2944 6556
rect 2944 6500 2948 6556
rect 2884 6496 2948 6500
rect 2964 6556 3028 6560
rect 2964 6500 2968 6556
rect 2968 6500 3024 6556
rect 3024 6500 3028 6556
rect 2964 6496 3028 6500
rect 3044 6556 3108 6560
rect 3044 6500 3048 6556
rect 3048 6500 3104 6556
rect 3104 6500 3108 6556
rect 3044 6496 3108 6500
rect 3124 6556 3188 6560
rect 3124 6500 3128 6556
rect 3128 6500 3184 6556
rect 3184 6500 3188 6556
rect 3124 6496 3188 6500
rect 4816 6556 4880 6560
rect 4816 6500 4820 6556
rect 4820 6500 4876 6556
rect 4876 6500 4880 6556
rect 4816 6496 4880 6500
rect 4896 6556 4960 6560
rect 4896 6500 4900 6556
rect 4900 6500 4956 6556
rect 4956 6500 4960 6556
rect 4896 6496 4960 6500
rect 4976 6556 5040 6560
rect 4976 6500 4980 6556
rect 4980 6500 5036 6556
rect 5036 6500 5040 6556
rect 4976 6496 5040 6500
rect 5056 6556 5120 6560
rect 5056 6500 5060 6556
rect 5060 6500 5116 6556
rect 5116 6500 5120 6556
rect 5056 6496 5120 6500
rect 6748 6556 6812 6560
rect 6748 6500 6752 6556
rect 6752 6500 6808 6556
rect 6808 6500 6812 6556
rect 6748 6496 6812 6500
rect 6828 6556 6892 6560
rect 6828 6500 6832 6556
rect 6832 6500 6888 6556
rect 6888 6500 6892 6556
rect 6828 6496 6892 6500
rect 6908 6556 6972 6560
rect 6908 6500 6912 6556
rect 6912 6500 6968 6556
rect 6968 6500 6972 6556
rect 6908 6496 6972 6500
rect 6988 6556 7052 6560
rect 6988 6500 6992 6556
rect 6992 6500 7048 6556
rect 7048 6500 7052 6556
rect 6988 6496 7052 6500
rect 8680 6556 8744 6560
rect 8680 6500 8684 6556
rect 8684 6500 8740 6556
rect 8740 6500 8744 6556
rect 8680 6496 8744 6500
rect 8760 6556 8824 6560
rect 8760 6500 8764 6556
rect 8764 6500 8820 6556
rect 8820 6500 8824 6556
rect 8760 6496 8824 6500
rect 8840 6556 8904 6560
rect 8840 6500 8844 6556
rect 8844 6500 8900 6556
rect 8900 6500 8904 6556
rect 8840 6496 8904 6500
rect 8920 6556 8984 6560
rect 8920 6500 8924 6556
rect 8924 6500 8980 6556
rect 8980 6500 8984 6556
rect 8920 6496 8984 6500
rect 1918 6012 1982 6016
rect 1918 5956 1922 6012
rect 1922 5956 1978 6012
rect 1978 5956 1982 6012
rect 1918 5952 1982 5956
rect 1998 6012 2062 6016
rect 1998 5956 2002 6012
rect 2002 5956 2058 6012
rect 2058 5956 2062 6012
rect 1998 5952 2062 5956
rect 2078 6012 2142 6016
rect 2078 5956 2082 6012
rect 2082 5956 2138 6012
rect 2138 5956 2142 6012
rect 2078 5952 2142 5956
rect 2158 6012 2222 6016
rect 2158 5956 2162 6012
rect 2162 5956 2218 6012
rect 2218 5956 2222 6012
rect 2158 5952 2222 5956
rect 3850 6012 3914 6016
rect 3850 5956 3854 6012
rect 3854 5956 3910 6012
rect 3910 5956 3914 6012
rect 3850 5952 3914 5956
rect 3930 6012 3994 6016
rect 3930 5956 3934 6012
rect 3934 5956 3990 6012
rect 3990 5956 3994 6012
rect 3930 5952 3994 5956
rect 4010 6012 4074 6016
rect 4010 5956 4014 6012
rect 4014 5956 4070 6012
rect 4070 5956 4074 6012
rect 4010 5952 4074 5956
rect 4090 6012 4154 6016
rect 4090 5956 4094 6012
rect 4094 5956 4150 6012
rect 4150 5956 4154 6012
rect 4090 5952 4154 5956
rect 5782 6012 5846 6016
rect 5782 5956 5786 6012
rect 5786 5956 5842 6012
rect 5842 5956 5846 6012
rect 5782 5952 5846 5956
rect 5862 6012 5926 6016
rect 5862 5956 5866 6012
rect 5866 5956 5922 6012
rect 5922 5956 5926 6012
rect 5862 5952 5926 5956
rect 5942 6012 6006 6016
rect 5942 5956 5946 6012
rect 5946 5956 6002 6012
rect 6002 5956 6006 6012
rect 5942 5952 6006 5956
rect 6022 6012 6086 6016
rect 6022 5956 6026 6012
rect 6026 5956 6082 6012
rect 6082 5956 6086 6012
rect 6022 5952 6086 5956
rect 7714 6012 7778 6016
rect 7714 5956 7718 6012
rect 7718 5956 7774 6012
rect 7774 5956 7778 6012
rect 7714 5952 7778 5956
rect 7794 6012 7858 6016
rect 7794 5956 7798 6012
rect 7798 5956 7854 6012
rect 7854 5956 7858 6012
rect 7794 5952 7858 5956
rect 7874 6012 7938 6016
rect 7874 5956 7878 6012
rect 7878 5956 7934 6012
rect 7934 5956 7938 6012
rect 7874 5952 7938 5956
rect 7954 6012 8018 6016
rect 7954 5956 7958 6012
rect 7958 5956 8014 6012
rect 8014 5956 8018 6012
rect 7954 5952 8018 5956
rect 2884 5468 2948 5472
rect 2884 5412 2888 5468
rect 2888 5412 2944 5468
rect 2944 5412 2948 5468
rect 2884 5408 2948 5412
rect 2964 5468 3028 5472
rect 2964 5412 2968 5468
rect 2968 5412 3024 5468
rect 3024 5412 3028 5468
rect 2964 5408 3028 5412
rect 3044 5468 3108 5472
rect 3044 5412 3048 5468
rect 3048 5412 3104 5468
rect 3104 5412 3108 5468
rect 3044 5408 3108 5412
rect 3124 5468 3188 5472
rect 3124 5412 3128 5468
rect 3128 5412 3184 5468
rect 3184 5412 3188 5468
rect 3124 5408 3188 5412
rect 4816 5468 4880 5472
rect 4816 5412 4820 5468
rect 4820 5412 4876 5468
rect 4876 5412 4880 5468
rect 4816 5408 4880 5412
rect 4896 5468 4960 5472
rect 4896 5412 4900 5468
rect 4900 5412 4956 5468
rect 4956 5412 4960 5468
rect 4896 5408 4960 5412
rect 4976 5468 5040 5472
rect 4976 5412 4980 5468
rect 4980 5412 5036 5468
rect 5036 5412 5040 5468
rect 4976 5408 5040 5412
rect 5056 5468 5120 5472
rect 5056 5412 5060 5468
rect 5060 5412 5116 5468
rect 5116 5412 5120 5468
rect 5056 5408 5120 5412
rect 6748 5468 6812 5472
rect 6748 5412 6752 5468
rect 6752 5412 6808 5468
rect 6808 5412 6812 5468
rect 6748 5408 6812 5412
rect 6828 5468 6892 5472
rect 6828 5412 6832 5468
rect 6832 5412 6888 5468
rect 6888 5412 6892 5468
rect 6828 5408 6892 5412
rect 6908 5468 6972 5472
rect 6908 5412 6912 5468
rect 6912 5412 6968 5468
rect 6968 5412 6972 5468
rect 6908 5408 6972 5412
rect 6988 5468 7052 5472
rect 6988 5412 6992 5468
rect 6992 5412 7048 5468
rect 7048 5412 7052 5468
rect 6988 5408 7052 5412
rect 8680 5468 8744 5472
rect 8680 5412 8684 5468
rect 8684 5412 8740 5468
rect 8740 5412 8744 5468
rect 8680 5408 8744 5412
rect 8760 5468 8824 5472
rect 8760 5412 8764 5468
rect 8764 5412 8820 5468
rect 8820 5412 8824 5468
rect 8760 5408 8824 5412
rect 8840 5468 8904 5472
rect 8840 5412 8844 5468
rect 8844 5412 8900 5468
rect 8900 5412 8904 5468
rect 8840 5408 8904 5412
rect 8920 5468 8984 5472
rect 8920 5412 8924 5468
rect 8924 5412 8980 5468
rect 8980 5412 8984 5468
rect 8920 5408 8984 5412
rect 1918 4924 1982 4928
rect 1918 4868 1922 4924
rect 1922 4868 1978 4924
rect 1978 4868 1982 4924
rect 1918 4864 1982 4868
rect 1998 4924 2062 4928
rect 1998 4868 2002 4924
rect 2002 4868 2058 4924
rect 2058 4868 2062 4924
rect 1998 4864 2062 4868
rect 2078 4924 2142 4928
rect 2078 4868 2082 4924
rect 2082 4868 2138 4924
rect 2138 4868 2142 4924
rect 2078 4864 2142 4868
rect 2158 4924 2222 4928
rect 2158 4868 2162 4924
rect 2162 4868 2218 4924
rect 2218 4868 2222 4924
rect 2158 4864 2222 4868
rect 3850 4924 3914 4928
rect 3850 4868 3854 4924
rect 3854 4868 3910 4924
rect 3910 4868 3914 4924
rect 3850 4864 3914 4868
rect 3930 4924 3994 4928
rect 3930 4868 3934 4924
rect 3934 4868 3990 4924
rect 3990 4868 3994 4924
rect 3930 4864 3994 4868
rect 4010 4924 4074 4928
rect 4010 4868 4014 4924
rect 4014 4868 4070 4924
rect 4070 4868 4074 4924
rect 4010 4864 4074 4868
rect 4090 4924 4154 4928
rect 4090 4868 4094 4924
rect 4094 4868 4150 4924
rect 4150 4868 4154 4924
rect 4090 4864 4154 4868
rect 5782 4924 5846 4928
rect 5782 4868 5786 4924
rect 5786 4868 5842 4924
rect 5842 4868 5846 4924
rect 5782 4864 5846 4868
rect 5862 4924 5926 4928
rect 5862 4868 5866 4924
rect 5866 4868 5922 4924
rect 5922 4868 5926 4924
rect 5862 4864 5926 4868
rect 5942 4924 6006 4928
rect 5942 4868 5946 4924
rect 5946 4868 6002 4924
rect 6002 4868 6006 4924
rect 5942 4864 6006 4868
rect 6022 4924 6086 4928
rect 6022 4868 6026 4924
rect 6026 4868 6082 4924
rect 6082 4868 6086 4924
rect 6022 4864 6086 4868
rect 7714 4924 7778 4928
rect 7714 4868 7718 4924
rect 7718 4868 7774 4924
rect 7774 4868 7778 4924
rect 7714 4864 7778 4868
rect 7794 4924 7858 4928
rect 7794 4868 7798 4924
rect 7798 4868 7854 4924
rect 7854 4868 7858 4924
rect 7794 4864 7858 4868
rect 7874 4924 7938 4928
rect 7874 4868 7878 4924
rect 7878 4868 7934 4924
rect 7934 4868 7938 4924
rect 7874 4864 7938 4868
rect 7954 4924 8018 4928
rect 7954 4868 7958 4924
rect 7958 4868 8014 4924
rect 8014 4868 8018 4924
rect 7954 4864 8018 4868
rect 2884 4380 2948 4384
rect 2884 4324 2888 4380
rect 2888 4324 2944 4380
rect 2944 4324 2948 4380
rect 2884 4320 2948 4324
rect 2964 4380 3028 4384
rect 2964 4324 2968 4380
rect 2968 4324 3024 4380
rect 3024 4324 3028 4380
rect 2964 4320 3028 4324
rect 3044 4380 3108 4384
rect 3044 4324 3048 4380
rect 3048 4324 3104 4380
rect 3104 4324 3108 4380
rect 3044 4320 3108 4324
rect 3124 4380 3188 4384
rect 3124 4324 3128 4380
rect 3128 4324 3184 4380
rect 3184 4324 3188 4380
rect 3124 4320 3188 4324
rect 4816 4380 4880 4384
rect 4816 4324 4820 4380
rect 4820 4324 4876 4380
rect 4876 4324 4880 4380
rect 4816 4320 4880 4324
rect 4896 4380 4960 4384
rect 4896 4324 4900 4380
rect 4900 4324 4956 4380
rect 4956 4324 4960 4380
rect 4896 4320 4960 4324
rect 4976 4380 5040 4384
rect 4976 4324 4980 4380
rect 4980 4324 5036 4380
rect 5036 4324 5040 4380
rect 4976 4320 5040 4324
rect 5056 4380 5120 4384
rect 5056 4324 5060 4380
rect 5060 4324 5116 4380
rect 5116 4324 5120 4380
rect 5056 4320 5120 4324
rect 6748 4380 6812 4384
rect 6748 4324 6752 4380
rect 6752 4324 6808 4380
rect 6808 4324 6812 4380
rect 6748 4320 6812 4324
rect 6828 4380 6892 4384
rect 6828 4324 6832 4380
rect 6832 4324 6888 4380
rect 6888 4324 6892 4380
rect 6828 4320 6892 4324
rect 6908 4380 6972 4384
rect 6908 4324 6912 4380
rect 6912 4324 6968 4380
rect 6968 4324 6972 4380
rect 6908 4320 6972 4324
rect 6988 4380 7052 4384
rect 6988 4324 6992 4380
rect 6992 4324 7048 4380
rect 7048 4324 7052 4380
rect 6988 4320 7052 4324
rect 8680 4380 8744 4384
rect 8680 4324 8684 4380
rect 8684 4324 8740 4380
rect 8740 4324 8744 4380
rect 8680 4320 8744 4324
rect 8760 4380 8824 4384
rect 8760 4324 8764 4380
rect 8764 4324 8820 4380
rect 8820 4324 8824 4380
rect 8760 4320 8824 4324
rect 8840 4380 8904 4384
rect 8840 4324 8844 4380
rect 8844 4324 8900 4380
rect 8900 4324 8904 4380
rect 8840 4320 8904 4324
rect 8920 4380 8984 4384
rect 8920 4324 8924 4380
rect 8924 4324 8980 4380
rect 8980 4324 8984 4380
rect 8920 4320 8984 4324
rect 1918 3836 1982 3840
rect 1918 3780 1922 3836
rect 1922 3780 1978 3836
rect 1978 3780 1982 3836
rect 1918 3776 1982 3780
rect 1998 3836 2062 3840
rect 1998 3780 2002 3836
rect 2002 3780 2058 3836
rect 2058 3780 2062 3836
rect 1998 3776 2062 3780
rect 2078 3836 2142 3840
rect 2078 3780 2082 3836
rect 2082 3780 2138 3836
rect 2138 3780 2142 3836
rect 2078 3776 2142 3780
rect 2158 3836 2222 3840
rect 2158 3780 2162 3836
rect 2162 3780 2218 3836
rect 2218 3780 2222 3836
rect 2158 3776 2222 3780
rect 3850 3836 3914 3840
rect 3850 3780 3854 3836
rect 3854 3780 3910 3836
rect 3910 3780 3914 3836
rect 3850 3776 3914 3780
rect 3930 3836 3994 3840
rect 3930 3780 3934 3836
rect 3934 3780 3990 3836
rect 3990 3780 3994 3836
rect 3930 3776 3994 3780
rect 4010 3836 4074 3840
rect 4010 3780 4014 3836
rect 4014 3780 4070 3836
rect 4070 3780 4074 3836
rect 4010 3776 4074 3780
rect 4090 3836 4154 3840
rect 4090 3780 4094 3836
rect 4094 3780 4150 3836
rect 4150 3780 4154 3836
rect 4090 3776 4154 3780
rect 5782 3836 5846 3840
rect 5782 3780 5786 3836
rect 5786 3780 5842 3836
rect 5842 3780 5846 3836
rect 5782 3776 5846 3780
rect 5862 3836 5926 3840
rect 5862 3780 5866 3836
rect 5866 3780 5922 3836
rect 5922 3780 5926 3836
rect 5862 3776 5926 3780
rect 5942 3836 6006 3840
rect 5942 3780 5946 3836
rect 5946 3780 6002 3836
rect 6002 3780 6006 3836
rect 5942 3776 6006 3780
rect 6022 3836 6086 3840
rect 6022 3780 6026 3836
rect 6026 3780 6082 3836
rect 6082 3780 6086 3836
rect 6022 3776 6086 3780
rect 7714 3836 7778 3840
rect 7714 3780 7718 3836
rect 7718 3780 7774 3836
rect 7774 3780 7778 3836
rect 7714 3776 7778 3780
rect 7794 3836 7858 3840
rect 7794 3780 7798 3836
rect 7798 3780 7854 3836
rect 7854 3780 7858 3836
rect 7794 3776 7858 3780
rect 7874 3836 7938 3840
rect 7874 3780 7878 3836
rect 7878 3780 7934 3836
rect 7934 3780 7938 3836
rect 7874 3776 7938 3780
rect 7954 3836 8018 3840
rect 7954 3780 7958 3836
rect 7958 3780 8014 3836
rect 8014 3780 8018 3836
rect 7954 3776 8018 3780
rect 2884 3292 2948 3296
rect 2884 3236 2888 3292
rect 2888 3236 2944 3292
rect 2944 3236 2948 3292
rect 2884 3232 2948 3236
rect 2964 3292 3028 3296
rect 2964 3236 2968 3292
rect 2968 3236 3024 3292
rect 3024 3236 3028 3292
rect 2964 3232 3028 3236
rect 3044 3292 3108 3296
rect 3044 3236 3048 3292
rect 3048 3236 3104 3292
rect 3104 3236 3108 3292
rect 3044 3232 3108 3236
rect 3124 3292 3188 3296
rect 3124 3236 3128 3292
rect 3128 3236 3184 3292
rect 3184 3236 3188 3292
rect 3124 3232 3188 3236
rect 4816 3292 4880 3296
rect 4816 3236 4820 3292
rect 4820 3236 4876 3292
rect 4876 3236 4880 3292
rect 4816 3232 4880 3236
rect 4896 3292 4960 3296
rect 4896 3236 4900 3292
rect 4900 3236 4956 3292
rect 4956 3236 4960 3292
rect 4896 3232 4960 3236
rect 4976 3292 5040 3296
rect 4976 3236 4980 3292
rect 4980 3236 5036 3292
rect 5036 3236 5040 3292
rect 4976 3232 5040 3236
rect 5056 3292 5120 3296
rect 5056 3236 5060 3292
rect 5060 3236 5116 3292
rect 5116 3236 5120 3292
rect 5056 3232 5120 3236
rect 6748 3292 6812 3296
rect 6748 3236 6752 3292
rect 6752 3236 6808 3292
rect 6808 3236 6812 3292
rect 6748 3232 6812 3236
rect 6828 3292 6892 3296
rect 6828 3236 6832 3292
rect 6832 3236 6888 3292
rect 6888 3236 6892 3292
rect 6828 3232 6892 3236
rect 6908 3292 6972 3296
rect 6908 3236 6912 3292
rect 6912 3236 6968 3292
rect 6968 3236 6972 3292
rect 6908 3232 6972 3236
rect 6988 3292 7052 3296
rect 6988 3236 6992 3292
rect 6992 3236 7048 3292
rect 7048 3236 7052 3292
rect 6988 3232 7052 3236
rect 8680 3292 8744 3296
rect 8680 3236 8684 3292
rect 8684 3236 8740 3292
rect 8740 3236 8744 3292
rect 8680 3232 8744 3236
rect 8760 3292 8824 3296
rect 8760 3236 8764 3292
rect 8764 3236 8820 3292
rect 8820 3236 8824 3292
rect 8760 3232 8824 3236
rect 8840 3292 8904 3296
rect 8840 3236 8844 3292
rect 8844 3236 8900 3292
rect 8900 3236 8904 3292
rect 8840 3232 8904 3236
rect 8920 3292 8984 3296
rect 8920 3236 8924 3292
rect 8924 3236 8980 3292
rect 8980 3236 8984 3292
rect 8920 3232 8984 3236
rect 1918 2748 1982 2752
rect 1918 2692 1922 2748
rect 1922 2692 1978 2748
rect 1978 2692 1982 2748
rect 1918 2688 1982 2692
rect 1998 2748 2062 2752
rect 1998 2692 2002 2748
rect 2002 2692 2058 2748
rect 2058 2692 2062 2748
rect 1998 2688 2062 2692
rect 2078 2748 2142 2752
rect 2078 2692 2082 2748
rect 2082 2692 2138 2748
rect 2138 2692 2142 2748
rect 2078 2688 2142 2692
rect 2158 2748 2222 2752
rect 2158 2692 2162 2748
rect 2162 2692 2218 2748
rect 2218 2692 2222 2748
rect 2158 2688 2222 2692
rect 3850 2748 3914 2752
rect 3850 2692 3854 2748
rect 3854 2692 3910 2748
rect 3910 2692 3914 2748
rect 3850 2688 3914 2692
rect 3930 2748 3994 2752
rect 3930 2692 3934 2748
rect 3934 2692 3990 2748
rect 3990 2692 3994 2748
rect 3930 2688 3994 2692
rect 4010 2748 4074 2752
rect 4010 2692 4014 2748
rect 4014 2692 4070 2748
rect 4070 2692 4074 2748
rect 4010 2688 4074 2692
rect 4090 2748 4154 2752
rect 4090 2692 4094 2748
rect 4094 2692 4150 2748
rect 4150 2692 4154 2748
rect 4090 2688 4154 2692
rect 5782 2748 5846 2752
rect 5782 2692 5786 2748
rect 5786 2692 5842 2748
rect 5842 2692 5846 2748
rect 5782 2688 5846 2692
rect 5862 2748 5926 2752
rect 5862 2692 5866 2748
rect 5866 2692 5922 2748
rect 5922 2692 5926 2748
rect 5862 2688 5926 2692
rect 5942 2748 6006 2752
rect 5942 2692 5946 2748
rect 5946 2692 6002 2748
rect 6002 2692 6006 2748
rect 5942 2688 6006 2692
rect 6022 2748 6086 2752
rect 6022 2692 6026 2748
rect 6026 2692 6082 2748
rect 6082 2692 6086 2748
rect 6022 2688 6086 2692
rect 7714 2748 7778 2752
rect 7714 2692 7718 2748
rect 7718 2692 7774 2748
rect 7774 2692 7778 2748
rect 7714 2688 7778 2692
rect 7794 2748 7858 2752
rect 7794 2692 7798 2748
rect 7798 2692 7854 2748
rect 7854 2692 7858 2748
rect 7794 2688 7858 2692
rect 7874 2748 7938 2752
rect 7874 2692 7878 2748
rect 7878 2692 7934 2748
rect 7934 2692 7938 2748
rect 7874 2688 7938 2692
rect 7954 2748 8018 2752
rect 7954 2692 7958 2748
rect 7958 2692 8014 2748
rect 8014 2692 8018 2748
rect 7954 2688 8018 2692
rect 2884 2204 2948 2208
rect 2884 2148 2888 2204
rect 2888 2148 2944 2204
rect 2944 2148 2948 2204
rect 2884 2144 2948 2148
rect 2964 2204 3028 2208
rect 2964 2148 2968 2204
rect 2968 2148 3024 2204
rect 3024 2148 3028 2204
rect 2964 2144 3028 2148
rect 3044 2204 3108 2208
rect 3044 2148 3048 2204
rect 3048 2148 3104 2204
rect 3104 2148 3108 2204
rect 3044 2144 3108 2148
rect 3124 2204 3188 2208
rect 3124 2148 3128 2204
rect 3128 2148 3184 2204
rect 3184 2148 3188 2204
rect 3124 2144 3188 2148
rect 4816 2204 4880 2208
rect 4816 2148 4820 2204
rect 4820 2148 4876 2204
rect 4876 2148 4880 2204
rect 4816 2144 4880 2148
rect 4896 2204 4960 2208
rect 4896 2148 4900 2204
rect 4900 2148 4956 2204
rect 4956 2148 4960 2204
rect 4896 2144 4960 2148
rect 4976 2204 5040 2208
rect 4976 2148 4980 2204
rect 4980 2148 5036 2204
rect 5036 2148 5040 2204
rect 4976 2144 5040 2148
rect 5056 2204 5120 2208
rect 5056 2148 5060 2204
rect 5060 2148 5116 2204
rect 5116 2148 5120 2204
rect 5056 2144 5120 2148
rect 6748 2204 6812 2208
rect 6748 2148 6752 2204
rect 6752 2148 6808 2204
rect 6808 2148 6812 2204
rect 6748 2144 6812 2148
rect 6828 2204 6892 2208
rect 6828 2148 6832 2204
rect 6832 2148 6888 2204
rect 6888 2148 6892 2204
rect 6828 2144 6892 2148
rect 6908 2204 6972 2208
rect 6908 2148 6912 2204
rect 6912 2148 6968 2204
rect 6968 2148 6972 2204
rect 6908 2144 6972 2148
rect 6988 2204 7052 2208
rect 6988 2148 6992 2204
rect 6992 2148 7048 2204
rect 7048 2148 7052 2204
rect 6988 2144 7052 2148
rect 8680 2204 8744 2208
rect 8680 2148 8684 2204
rect 8684 2148 8740 2204
rect 8740 2148 8744 2204
rect 8680 2144 8744 2148
rect 8760 2204 8824 2208
rect 8760 2148 8764 2204
rect 8764 2148 8820 2204
rect 8820 2148 8824 2204
rect 8760 2144 8824 2148
rect 8840 2204 8904 2208
rect 8840 2148 8844 2204
rect 8844 2148 8900 2204
rect 8900 2148 8904 2204
rect 8840 2144 8904 2148
rect 8920 2204 8984 2208
rect 8920 2148 8924 2204
rect 8924 2148 8980 2204
rect 8980 2148 8984 2204
rect 8920 2144 8984 2148
<< metal4 >>
rect 1910 7104 2230 7664
rect 1910 7040 1918 7104
rect 1982 7040 1998 7104
rect 2062 7040 2078 7104
rect 2142 7040 2158 7104
rect 2222 7040 2230 7104
rect 1910 6016 2230 7040
rect 1910 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2230 6016
rect 1910 4928 2230 5952
rect 1910 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2230 4928
rect 1910 3840 2230 4864
rect 1910 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2230 3840
rect 1910 2752 2230 3776
rect 1910 2688 1918 2752
rect 1982 2688 1998 2752
rect 2062 2688 2078 2752
rect 2142 2688 2158 2752
rect 2222 2688 2230 2752
rect 1910 2128 2230 2688
rect 2876 7648 3196 7664
rect 2876 7584 2884 7648
rect 2948 7584 2964 7648
rect 3028 7584 3044 7648
rect 3108 7584 3124 7648
rect 3188 7584 3196 7648
rect 2876 6560 3196 7584
rect 2876 6496 2884 6560
rect 2948 6496 2964 6560
rect 3028 6496 3044 6560
rect 3108 6496 3124 6560
rect 3188 6496 3196 6560
rect 2876 5472 3196 6496
rect 2876 5408 2884 5472
rect 2948 5408 2964 5472
rect 3028 5408 3044 5472
rect 3108 5408 3124 5472
rect 3188 5408 3196 5472
rect 2876 4384 3196 5408
rect 2876 4320 2884 4384
rect 2948 4320 2964 4384
rect 3028 4320 3044 4384
rect 3108 4320 3124 4384
rect 3188 4320 3196 4384
rect 2876 3296 3196 4320
rect 2876 3232 2884 3296
rect 2948 3232 2964 3296
rect 3028 3232 3044 3296
rect 3108 3232 3124 3296
rect 3188 3232 3196 3296
rect 2876 2208 3196 3232
rect 2876 2144 2884 2208
rect 2948 2144 2964 2208
rect 3028 2144 3044 2208
rect 3108 2144 3124 2208
rect 3188 2144 3196 2208
rect 2876 2128 3196 2144
rect 3842 7104 4162 7664
rect 3842 7040 3850 7104
rect 3914 7040 3930 7104
rect 3994 7040 4010 7104
rect 4074 7040 4090 7104
rect 4154 7040 4162 7104
rect 3842 6016 4162 7040
rect 3842 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4162 6016
rect 3842 4928 4162 5952
rect 3842 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4162 4928
rect 3842 3840 4162 4864
rect 3842 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4162 3840
rect 3842 2752 4162 3776
rect 3842 2688 3850 2752
rect 3914 2688 3930 2752
rect 3994 2688 4010 2752
rect 4074 2688 4090 2752
rect 4154 2688 4162 2752
rect 3842 2128 4162 2688
rect 4808 7648 5128 7664
rect 4808 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5128 7648
rect 4808 6560 5128 7584
rect 4808 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5128 6560
rect 4808 5472 5128 6496
rect 4808 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5128 5472
rect 4808 4384 5128 5408
rect 4808 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5128 4384
rect 4808 3296 5128 4320
rect 4808 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5128 3296
rect 4808 2208 5128 3232
rect 4808 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5128 2208
rect 4808 2128 5128 2144
rect 5774 7104 6094 7664
rect 5774 7040 5782 7104
rect 5846 7040 5862 7104
rect 5926 7040 5942 7104
rect 6006 7040 6022 7104
rect 6086 7040 6094 7104
rect 5774 6016 6094 7040
rect 5774 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6094 6016
rect 5774 4928 6094 5952
rect 5774 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6094 4928
rect 5774 3840 6094 4864
rect 5774 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6094 3840
rect 5774 2752 6094 3776
rect 5774 2688 5782 2752
rect 5846 2688 5862 2752
rect 5926 2688 5942 2752
rect 6006 2688 6022 2752
rect 6086 2688 6094 2752
rect 5774 2128 6094 2688
rect 6740 7648 7060 7664
rect 6740 7584 6748 7648
rect 6812 7584 6828 7648
rect 6892 7584 6908 7648
rect 6972 7584 6988 7648
rect 7052 7584 7060 7648
rect 6740 6560 7060 7584
rect 6740 6496 6748 6560
rect 6812 6496 6828 6560
rect 6892 6496 6908 6560
rect 6972 6496 6988 6560
rect 7052 6496 7060 6560
rect 6740 5472 7060 6496
rect 6740 5408 6748 5472
rect 6812 5408 6828 5472
rect 6892 5408 6908 5472
rect 6972 5408 6988 5472
rect 7052 5408 7060 5472
rect 6740 4384 7060 5408
rect 6740 4320 6748 4384
rect 6812 4320 6828 4384
rect 6892 4320 6908 4384
rect 6972 4320 6988 4384
rect 7052 4320 7060 4384
rect 6740 3296 7060 4320
rect 6740 3232 6748 3296
rect 6812 3232 6828 3296
rect 6892 3232 6908 3296
rect 6972 3232 6988 3296
rect 7052 3232 7060 3296
rect 6740 2208 7060 3232
rect 6740 2144 6748 2208
rect 6812 2144 6828 2208
rect 6892 2144 6908 2208
rect 6972 2144 6988 2208
rect 7052 2144 7060 2208
rect 6740 2128 7060 2144
rect 7706 7104 8026 7664
rect 7706 7040 7714 7104
rect 7778 7040 7794 7104
rect 7858 7040 7874 7104
rect 7938 7040 7954 7104
rect 8018 7040 8026 7104
rect 7706 6016 8026 7040
rect 7706 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8026 6016
rect 7706 4928 8026 5952
rect 7706 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8026 4928
rect 7706 3840 8026 4864
rect 7706 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8026 3840
rect 7706 2752 8026 3776
rect 7706 2688 7714 2752
rect 7778 2688 7794 2752
rect 7858 2688 7874 2752
rect 7938 2688 7954 2752
rect 8018 2688 8026 2752
rect 7706 2128 8026 2688
rect 8672 7648 8992 7664
rect 8672 7584 8680 7648
rect 8744 7584 8760 7648
rect 8824 7584 8840 7648
rect 8904 7584 8920 7648
rect 8984 7584 8992 7648
rect 8672 6560 8992 7584
rect 8672 6496 8680 6560
rect 8744 6496 8760 6560
rect 8824 6496 8840 6560
rect 8904 6496 8920 6560
rect 8984 6496 8992 6560
rect 8672 5472 8992 6496
rect 8672 5408 8680 5472
rect 8744 5408 8760 5472
rect 8824 5408 8840 5472
rect 8904 5408 8920 5472
rect 8984 5408 8992 5472
rect 8672 4384 8992 5408
rect 8672 4320 8680 4384
rect 8744 4320 8760 4384
rect 8824 4320 8840 4384
rect 8904 4320 8920 4384
rect 8984 4320 8992 4384
rect 8672 3296 8992 4320
rect 8672 3232 8680 3296
rect 8744 3232 8760 3296
rect 8824 3232 8840 3296
rect 8904 3232 8920 3296
rect 8984 3232 8992 3296
rect 8672 2208 8992 3232
rect 8672 2144 8680 2208
rect 8744 2144 8760 2208
rect 8824 2144 8840 2208
rect 8904 2144 8920 2208
rect 8984 2144 8992 2208
rect 8672 2128 8992 2144
use sky130_fd_sc_hd__inv_2  _08_
timestamp 0
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _09_
timestamp 0
transform -1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _10_
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _11_
timestamp 0
transform 1 0 3864 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _12_
timestamp 0
transform 1 0 5336 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _13_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _14_
timestamp 0
transform -1 0 5336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _15_
timestamp 0
transform -1 0 5520 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _16_
timestamp 0
transform 1 0 6532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _17_
timestamp 0
transform 1 0 3772 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _18_
timestamp 0
transform -1 0 5244 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 4692 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 6716 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 0
transform -1 0 7268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_11
timestamp 0
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_45
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_57
timestamp 0
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_69
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_45
timestamp 0
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 0
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_75
timestamp 0
transform 1 0 8004 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_59
timestamp 0
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_67
timestamp 0
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_79
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_21
timestamp 0
transform 1 0 3036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_26
timestamp 0
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 0
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_46
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 0
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_65
timestamp 0
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform -1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 754 9200 810 10000 0 FreeSans 280 90 0 0 D[0]
port 1 nsew
flabel metal2 s 1950 9200 2006 10000 0 FreeSans 280 90 0 0 D[1]
port 2 nsew
flabel metal2 s 3146 9200 3202 10000 0 FreeSans 280 90 0 0 D[2]
port 3 nsew
flabel metal2 s 4342 9200 4398 10000 0 FreeSans 280 90 0 0 D[3]
port 4 nsew
flabel metal2 s 5538 9200 5594 10000 0 FreeSans 280 90 0 0 D[4]
port 5 nsew
flabel metal2 s 6734 9200 6790 10000 0 FreeSans 280 90 0 0 D[5]
port 6 nsew
flabel metal2 s 7930 9200 7986 10000 0 FreeSans 280 90 0 0 D[6]
port 7 nsew
flabel metal2 s 9126 9200 9182 10000 0 FreeSans 280 90 0 0 D[7]
port 8 nsew
flabel metal2 s 1674 0 1730 800 0 FreeSans 280 90 0 0 O[0]
port 9 nsew
flabel metal2 s 4986 0 5042 800 0 FreeSans 280 90 0 0 O[1]
port 10 nsew
flabel metal2 s 8298 0 8354 800 0 FreeSans 280 90 0 0 O[2]
port 11 nsew
flabel metal4 s 8672 2128 8992 7664 0 FreeSans 2400 90 0 0 VGND
port 12 nsew
flabel metal4 s 6740 2128 7060 7664 0 FreeSans 2400 90 0 0 VGND
port 12 nsew
flabel metal4 s 4808 2128 5128 7664 0 FreeSans 2400 90 0 0 VGND
port 12 nsew
flabel metal4 s 2876 2128 3196 7664 0 FreeSans 2400 90 0 0 VGND
port 12 nsew
flabel metal4 s 7706 2128 8026 7664 0 FreeSans 2400 90 0 0 VPWR
port 13 nsew
flabel metal4 s 5774 2128 6094 7664 0 FreeSans 2400 90 0 0 VPWR
port 13 nsew
flabel metal4 s 3842 2128 4162 7664 0 FreeSans 2400 90 0 0 VPWR
port 13 nsew
flabel metal4 s 1910 2128 2230 7664 0 FreeSans 2400 90 0 0 VPWR
port 13 nsew
flabel metal3 s 0 4904 800 5024 0 FreeSans 600 0 0 0 clk
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1730901468
<< nwell >>
rect 1066 2159 8870 7633
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 1104 2128 9186 7664
<< metal2 >>
rect 754 9200 810 10000
rect 1950 9200 2006 10000
rect 3146 9200 3202 10000
rect 4342 9200 4398 10000
rect 5538 9200 5594 10000
rect 6734 9200 6790 10000
rect 7930 9200 7986 10000
rect 9126 9200 9182 10000
rect 1674 0 1730 800
rect 4986 0 5042 800
rect 8298 0 8354 800
<< obsm2 >>
rect 1676 9144 1894 9330
rect 2062 9144 3090 9330
rect 3258 9144 4286 9330
rect 4454 9144 5482 9330
rect 5650 9144 6678 9330
rect 6846 9144 7874 9330
rect 8042 9144 9070 9330
rect 1676 856 9180 9144
rect 1786 800 4930 856
rect 5098 800 8242 856
rect 8410 800 9180 856
<< metal3 >>
rect 0 4904 800 5024
<< obsm3 >>
rect 800 5104 8990 7649
rect 880 4824 8990 5104
rect 800 2143 8990 4824
<< metal4 >>
rect 1910 2128 2230 7664
rect 2876 2128 3196 7664
rect 3842 2128 4162 7664
rect 4808 2128 5128 7664
rect 5774 2128 6094 7664
rect 6740 2128 7060 7664
rect 7706 2128 8026 7664
rect 8672 2128 8992 7664
<< labels >>
rlabel metal2 s 754 9200 810 10000 6 D[0]
port 1 nsew signal input
rlabel metal2 s 1950 9200 2006 10000 6 D[1]
port 2 nsew signal input
rlabel metal2 s 3146 9200 3202 10000 6 D[2]
port 3 nsew signal input
rlabel metal2 s 4342 9200 4398 10000 6 D[3]
port 4 nsew signal input
rlabel metal2 s 5538 9200 5594 10000 6 D[4]
port 5 nsew signal input
rlabel metal2 s 6734 9200 6790 10000 6 D[5]
port 6 nsew signal input
rlabel metal2 s 7930 9200 7986 10000 6 D[6]
port 7 nsew signal input
rlabel metal2 s 9126 9200 9182 10000 6 D[7]
port 8 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 O[0]
port 9 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 O[1]
port 10 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 O[2]
port 11 nsew signal output
rlabel metal4 s 2876 2128 3196 7664 6 VGND
port 12 nsew ground bidirectional
rlabel metal4 s 4808 2128 5128 7664 6 VGND
port 12 nsew ground bidirectional
rlabel metal4 s 6740 2128 7060 7664 6 VGND
port 12 nsew ground bidirectional
rlabel metal4 s 8672 2128 8992 7664 6 VGND
port 12 nsew ground bidirectional
rlabel metal4 s 1910 2128 2230 7664 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 3842 2128 4162 7664 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 5774 2128 6094 7664 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 7706 2128 8026 7664 6 VPWR
port 13 nsew power bidirectional
rlabel metal3 s 0 4904 800 5024 6 clk
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 197646
string GDS_FILE /openlane/designs/priority_encoder/runs/RUN_2024.11.06_13.57.03/results/signoff/priority_encoder.magic.gds
string GDS_START 103356
<< end >>

